module reg8000 ( in, clk, rst, out );
	input[31:0] in;
	input clk;
	input rst;
	output[31:0] out;

	wire [31:0] r0_out;
	wire [31:0] r1_out;
	wire [31:0] r2_out;
	wire [31:0] r3_out;
	wire [31:0] r4_out;
	wire [31:0] r5_out;
	wire [31:0] r6_out;
	wire [31:0] r7_out;
	wire [31:0] r8_out;
	wire [31:0] r9_out;
	wire [31:0] r10_out;
	wire [31:0] r11_out;
	wire [31:0] r12_out;
	wire [31:0] r13_out;
	wire [31:0] r14_out;
	wire [31:0] r15_out;
	wire [31:0] r16_out;
	wire [31:0] r17_out;
	wire [31:0] r18_out;
	wire [31:0] r19_out;
	wire [31:0] r20_out;
	wire [31:0] r21_out;
	wire [31:0] r22_out;
	wire [31:0] r23_out;
	wire [31:0] r24_out;
	wire [31:0] r25_out;
	wire [31:0] r26_out;
	wire [31:0] r27_out;
	wire [31:0] r28_out;
	wire [31:0] r29_out;
	wire [31:0] r30_out;
	wire [31:0] r31_out;
	wire [31:0] r32_out;
	wire [31:0] r33_out;
	wire [31:0] r34_out;
	wire [31:0] r35_out;
	wire [31:0] r36_out;
	wire [31:0] r37_out;
	wire [31:0] r38_out;
	wire [31:0] r39_out;
	wire [31:0] r40_out;
	wire [31:0] r41_out;
	wire [31:0] r42_out;
	wire [31:0] r43_out;
	wire [31:0] r44_out;
	wire [31:0] r45_out;
	wire [31:0] r46_out;
	wire [31:0] r47_out;
	wire [31:0] r48_out;
	wire [31:0] r49_out;
	wire [31:0] r50_out;
	wire [31:0] r51_out;
	wire [31:0] r52_out;
	wire [31:0] r53_out;
	wire [31:0] r54_out;
	wire [31:0] r55_out;
	wire [31:0] r56_out;
	wire [31:0] r57_out;
	wire [31:0] r58_out;
	wire [31:0] r59_out;
	wire [31:0] r60_out;
	wire [31:0] r61_out;
	wire [31:0] r62_out;
	wire [31:0] r63_out;
	wire [31:0] r64_out;
	wire [31:0] r65_out;
	wire [31:0] r66_out;
	wire [31:0] r67_out;
	wire [31:0] r68_out;
	wire [31:0] r69_out;
	wire [31:0] r70_out;
	wire [31:0] r71_out;
	wire [31:0] r72_out;
	wire [31:0] r73_out;
	wire [31:0] r74_out;
	wire [31:0] r75_out;
	wire [31:0] r76_out;
	wire [31:0] r77_out;
	wire [31:0] r78_out;
	wire [31:0] r79_out;
	wire [31:0] r80_out;
	wire [31:0] r81_out;
	wire [31:0] r82_out;
	wire [31:0] r83_out;
	wire [31:0] r84_out;
	wire [31:0] r85_out;
	wire [31:0] r86_out;
	wire [31:0] r87_out;
	wire [31:0] r88_out;
	wire [31:0] r89_out;
	wire [31:0] r90_out;
	wire [31:0] r91_out;
	wire [31:0] r92_out;
	wire [31:0] r93_out;
	wire [31:0] r94_out;
	wire [31:0] r95_out;
	wire [31:0] r96_out;
	wire [31:0] r97_out;
	wire [31:0] r98_out;
	wire [31:0] r99_out;
	wire [31:0] r100_out;
	wire [31:0] r101_out;
	wire [31:0] r102_out;
	wire [31:0] r103_out;
	wire [31:0] r104_out;
	wire [31:0] r105_out;
	wire [31:0] r106_out;
	wire [31:0] r107_out;
	wire [31:0] r108_out;
	wire [31:0] r109_out;
	wire [31:0] r110_out;
	wire [31:0] r111_out;
	wire [31:0] r112_out;
	wire [31:0] r113_out;
	wire [31:0] r114_out;
	wire [31:0] r115_out;
	wire [31:0] r116_out;
	wire [31:0] r117_out;
	wire [31:0] r118_out;
	wire [31:0] r119_out;
	wire [31:0] r120_out;
	wire [31:0] r121_out;
	wire [31:0] r122_out;
	wire [31:0] r123_out;
	wire [31:0] r124_out;
	wire [31:0] r125_out;
	wire [31:0] r126_out;
	wire [31:0] r127_out;
	wire [31:0] r128_out;
	wire [31:0] r129_out;
	wire [31:0] r130_out;
	wire [31:0] r131_out;
	wire [31:0] r132_out;
	wire [31:0] r133_out;
	wire [31:0] r134_out;
	wire [31:0] r135_out;
	wire [31:0] r136_out;
	wire [31:0] r137_out;
	wire [31:0] r138_out;
	wire [31:0] r139_out;
	wire [31:0] r140_out;
	wire [31:0] r141_out;
	wire [31:0] r142_out;
	wire [31:0] r143_out;
	wire [31:0] r144_out;
	wire [31:0] r145_out;
	wire [31:0] r146_out;
	wire [31:0] r147_out;
	wire [31:0] r148_out;
	wire [31:0] r149_out;
	wire [31:0] r150_out;
	wire [31:0] r151_out;
	wire [31:0] r152_out;
	wire [31:0] r153_out;
	wire [31:0] r154_out;
	wire [31:0] r155_out;
	wire [31:0] r156_out;
	wire [31:0] r157_out;
	wire [31:0] r158_out;
	wire [31:0] r159_out;
	wire [31:0] r160_out;
	wire [31:0] r161_out;
	wire [31:0] r162_out;
	wire [31:0] r163_out;
	wire [31:0] r164_out;
	wire [31:0] r165_out;
	wire [31:0] r166_out;
	wire [31:0] r167_out;
	wire [31:0] r168_out;
	wire [31:0] r169_out;
	wire [31:0] r170_out;
	wire [31:0] r171_out;
	wire [31:0] r172_out;
	wire [31:0] r173_out;
	wire [31:0] r174_out;
	wire [31:0] r175_out;
	wire [31:0] r176_out;
	wire [31:0] r177_out;
	wire [31:0] r178_out;
	wire [31:0] r179_out;
	wire [31:0] r180_out;
	wire [31:0] r181_out;
	wire [31:0] r182_out;
	wire [31:0] r183_out;
	wire [31:0] r184_out;
	wire [31:0] r185_out;
	wire [31:0] r186_out;
	wire [31:0] r187_out;
	wire [31:0] r188_out;
	wire [31:0] r189_out;
	wire [31:0] r190_out;
	wire [31:0] r191_out;
	wire [31:0] r192_out;
	wire [31:0] r193_out;
	wire [31:0] r194_out;
	wire [31:0] r195_out;
	wire [31:0] r196_out;
	wire [31:0] r197_out;
	wire [31:0] r198_out;
	wire [31:0] r199_out;
	wire [31:0] r200_out;
	wire [31:0] r201_out;
	wire [31:0] r202_out;
	wire [31:0] r203_out;
	wire [31:0] r204_out;
	wire [31:0] r205_out;
	wire [31:0] r206_out;
	wire [31:0] r207_out;
	wire [31:0] r208_out;
	wire [31:0] r209_out;
	wire [31:0] r210_out;
	wire [31:0] r211_out;
	wire [31:0] r212_out;
	wire [31:0] r213_out;
	wire [31:0] r214_out;
	wire [31:0] r215_out;
	wire [31:0] r216_out;
	wire [31:0] r217_out;
	wire [31:0] r218_out;
	wire [31:0] r219_out;
	wire [31:0] r220_out;
	wire [31:0] r221_out;
	wire [31:0] r222_out;
	wire [31:0] r223_out;
	wire [31:0] r224_out;
	wire [31:0] r225_out;
	wire [31:0] r226_out;
	wire [31:0] r227_out;
	wire [31:0] r228_out;
	wire [31:0] r229_out;
	wire [31:0] r230_out;
	wire [31:0] r231_out;
	wire [31:0] r232_out;
	wire [31:0] r233_out;
	wire [31:0] r234_out;
	wire [31:0] r235_out;
	wire [31:0] r236_out;
	wire [31:0] r237_out;
	wire [31:0] r238_out;
	wire [31:0] r239_out;
	wire [31:0] r240_out;
	wire [31:0] r241_out;
	wire [31:0] r242_out;
	wire [31:0] r243_out;
	wire [31:0] r244_out;
	wire [31:0] r245_out;
	wire [31:0] r246_out;
	wire [31:0] r247_out;
	wire [31:0] r248_out;
	wire [31:0] r249_out;
	wire [31:0] r250_out;
	wire [31:0] r251_out;
	wire [31:0] r252_out;
	wire [31:0] r253_out;
	wire [31:0] r254_out;
	wire [31:0] r255_out;
	wire [31:0] r256_out;
	wire [31:0] r257_out;
	wire [31:0] r258_out;
	wire [31:0] r259_out;
	wire [31:0] r260_out;
	wire [31:0] r261_out;
	wire [31:0] r262_out;
	wire [31:0] r263_out;
	wire [31:0] r264_out;
	wire [31:0] r265_out;
	wire [31:0] r266_out;
	wire [31:0] r267_out;
	wire [31:0] r268_out;
	wire [31:0] r269_out;
	wire [31:0] r270_out;
	wire [31:0] r271_out;
	wire [31:0] r272_out;
	wire [31:0] r273_out;
	wire [31:0] r274_out;
	wire [31:0] r275_out;
	wire [31:0] r276_out;
	wire [31:0] r277_out;
	wire [31:0] r278_out;
	wire [31:0] r279_out;
	wire [31:0] r280_out;
	wire [31:0] r281_out;
	wire [31:0] r282_out;
	wire [31:0] r283_out;
	wire [31:0] r284_out;
	wire [31:0] r285_out;
	wire [31:0] r286_out;
	wire [31:0] r287_out;
	wire [31:0] r288_out;
	wire [31:0] r289_out;
	wire [31:0] r290_out;
	wire [31:0] r291_out;
	wire [31:0] r292_out;
	wire [31:0] r293_out;
	wire [31:0] r294_out;
	wire [31:0] r295_out;
	wire [31:0] r296_out;
	wire [31:0] r297_out;
	wire [31:0] r298_out;
	wire [31:0] r299_out;
	wire [31:0] r300_out;
	wire [31:0] r301_out;
	wire [31:0] r302_out;
	wire [31:0] r303_out;
	wire [31:0] r304_out;
	wire [31:0] r305_out;
	wire [31:0] r306_out;
	wire [31:0] r307_out;
	wire [31:0] r308_out;
	wire [31:0] r309_out;
	wire [31:0] r310_out;
	wire [31:0] r311_out;
	wire [31:0] r312_out;
	wire [31:0] r313_out;
	wire [31:0] r314_out;
	wire [31:0] r315_out;
	wire [31:0] r316_out;
	wire [31:0] r317_out;
	wire [31:0] r318_out;
	wire [31:0] r319_out;
	wire [31:0] r320_out;
	wire [31:0] r321_out;
	wire [31:0] r322_out;
	wire [31:0] r323_out;
	wire [31:0] r324_out;
	wire [31:0] r325_out;
	wire [31:0] r326_out;
	wire [31:0] r327_out;
	wire [31:0] r328_out;
	wire [31:0] r329_out;
	wire [31:0] r330_out;
	wire [31:0] r331_out;
	wire [31:0] r332_out;
	wire [31:0] r333_out;
	wire [31:0] r334_out;
	wire [31:0] r335_out;
	wire [31:0] r336_out;
	wire [31:0] r337_out;
	wire [31:0] r338_out;
	wire [31:0] r339_out;
	wire [31:0] r340_out;
	wire [31:0] r341_out;
	wire [31:0] r342_out;
	wire [31:0] r343_out;
	wire [31:0] r344_out;
	wire [31:0] r345_out;
	wire [31:0] r346_out;
	wire [31:0] r347_out;
	wire [31:0] r348_out;
	wire [31:0] r349_out;
	wire [31:0] r350_out;
	wire [31:0] r351_out;
	wire [31:0] r352_out;
	wire [31:0] r353_out;
	wire [31:0] r354_out;
	wire [31:0] r355_out;
	wire [31:0] r356_out;
	wire [31:0] r357_out;
	wire [31:0] r358_out;
	wire [31:0] r359_out;
	wire [31:0] r360_out;
	wire [31:0] r361_out;
	wire [31:0] r362_out;
	wire [31:0] r363_out;
	wire [31:0] r364_out;
	wire [31:0] r365_out;
	wire [31:0] r366_out;
	wire [31:0] r367_out;
	wire [31:0] r368_out;
	wire [31:0] r369_out;
	wire [31:0] r370_out;
	wire [31:0] r371_out;
	wire [31:0] r372_out;
	wire [31:0] r373_out;
	wire [31:0] r374_out;
	wire [31:0] r375_out;
	wire [31:0] r376_out;
	wire [31:0] r377_out;
	wire [31:0] r378_out;
	wire [31:0] r379_out;
	wire [31:0] r380_out;
	wire [31:0] r381_out;
	wire [31:0] r382_out;
	wire [31:0] r383_out;
	wire [31:0] r384_out;
	wire [31:0] r385_out;
	wire [31:0] r386_out;
	wire [31:0] r387_out;
	wire [31:0] r388_out;
	wire [31:0] r389_out;
	wire [31:0] r390_out;
	wire [31:0] r391_out;
	wire [31:0] r392_out;
	wire [31:0] r393_out;
	wire [31:0] r394_out;
	wire [31:0] r395_out;
	wire [31:0] r396_out;
	wire [31:0] r397_out;
	wire [31:0] r398_out;
	wire [31:0] r399_out;
	wire [31:0] r400_out;
	wire [31:0] r401_out;
	wire [31:0] r402_out;
	wire [31:0] r403_out;
	wire [31:0] r404_out;
	wire [31:0] r405_out;
	wire [31:0] r406_out;
	wire [31:0] r407_out;
	wire [31:0] r408_out;
	wire [31:0] r409_out;
	wire [31:0] r410_out;
	wire [31:0] r411_out;
	wire [31:0] r412_out;
	wire [31:0] r413_out;
	wire [31:0] r414_out;
	wire [31:0] r415_out;
	wire [31:0] r416_out;
	wire [31:0] r417_out;
	wire [31:0] r418_out;
	wire [31:0] r419_out;
	wire [31:0] r420_out;
	wire [31:0] r421_out;
	wire [31:0] r422_out;
	wire [31:0] r423_out;
	wire [31:0] r424_out;
	wire [31:0] r425_out;
	wire [31:0] r426_out;
	wire [31:0] r427_out;
	wire [31:0] r428_out;
	wire [31:0] r429_out;
	wire [31:0] r430_out;
	wire [31:0] r431_out;
	wire [31:0] r432_out;
	wire [31:0] r433_out;
	wire [31:0] r434_out;
	wire [31:0] r435_out;
	wire [31:0] r436_out;
	wire [31:0] r437_out;
	wire [31:0] r438_out;
	wire [31:0] r439_out;
	wire [31:0] r440_out;
	wire [31:0] r441_out;
	wire [31:0] r442_out;
	wire [31:0] r443_out;
	wire [31:0] r444_out;
	wire [31:0] r445_out;
	wire [31:0] r446_out;
	wire [31:0] r447_out;
	wire [31:0] r448_out;
	wire [31:0] r449_out;
	wire [31:0] r450_out;
	wire [31:0] r451_out;
	wire [31:0] r452_out;
	wire [31:0] r453_out;
	wire [31:0] r454_out;
	wire [31:0] r455_out;
	wire [31:0] r456_out;
	wire [31:0] r457_out;
	wire [31:0] r458_out;
	wire [31:0] r459_out;
	wire [31:0] r460_out;
	wire [31:0] r461_out;
	wire [31:0] r462_out;
	wire [31:0] r463_out;
	wire [31:0] r464_out;
	wire [31:0] r465_out;
	wire [31:0] r466_out;
	wire [31:0] r467_out;
	wire [31:0] r468_out;
	wire [31:0] r469_out;
	wire [31:0] r470_out;
	wire [31:0] r471_out;
	wire [31:0] r472_out;
	wire [31:0] r473_out;
	wire [31:0] r474_out;
	wire [31:0] r475_out;
	wire [31:0] r476_out;
	wire [31:0] r477_out;
	wire [31:0] r478_out;
	wire [31:0] r479_out;
	wire [31:0] r480_out;
	wire [31:0] r481_out;
	wire [31:0] r482_out;
	wire [31:0] r483_out;
	wire [31:0] r484_out;
	wire [31:0] r485_out;
	wire [31:0] r486_out;
	wire [31:0] r487_out;
	wire [31:0] r488_out;
	wire [31:0] r489_out;
	wire [31:0] r490_out;
	wire [31:0] r491_out;
	wire [31:0] r492_out;
	wire [31:0] r493_out;
	wire [31:0] r494_out;
	wire [31:0] r495_out;
	wire [31:0] r496_out;
	wire [31:0] r497_out;
	wire [31:0] r498_out;
	wire [31:0] r499_out;
	wire [31:0] r500_out;
	wire [31:0] r501_out;
	wire [31:0] r502_out;
	wire [31:0] r503_out;
	wire [31:0] r504_out;
	wire [31:0] r505_out;
	wire [31:0] r506_out;
	wire [31:0] r507_out;
	wire [31:0] r508_out;
	wire [31:0] r509_out;
	wire [31:0] r510_out;
	wire [31:0] r511_out;
	wire [31:0] r512_out;
	wire [31:0] r513_out;
	wire [31:0] r514_out;
	wire [31:0] r515_out;
	wire [31:0] r516_out;
	wire [31:0] r517_out;
	wire [31:0] r518_out;
	wire [31:0] r519_out;
	wire [31:0] r520_out;
	wire [31:0] r521_out;
	wire [31:0] r522_out;
	wire [31:0] r523_out;
	wire [31:0] r524_out;
	wire [31:0] r525_out;
	wire [31:0] r526_out;
	wire [31:0] r527_out;
	wire [31:0] r528_out;
	wire [31:0] r529_out;
	wire [31:0] r530_out;
	wire [31:0] r531_out;
	wire [31:0] r532_out;
	wire [31:0] r533_out;
	wire [31:0] r534_out;
	wire [31:0] r535_out;
	wire [31:0] r536_out;
	wire [31:0] r537_out;
	wire [31:0] r538_out;
	wire [31:0] r539_out;
	wire [31:0] r540_out;
	wire [31:0] r541_out;
	wire [31:0] r542_out;
	wire [31:0] r543_out;
	wire [31:0] r544_out;
	wire [31:0] r545_out;
	wire [31:0] r546_out;
	wire [31:0] r547_out;
	wire [31:0] r548_out;
	wire [31:0] r549_out;
	wire [31:0] r550_out;
	wire [31:0] r551_out;
	wire [31:0] r552_out;
	wire [31:0] r553_out;
	wire [31:0] r554_out;
	wire [31:0] r555_out;
	wire [31:0] r556_out;
	wire [31:0] r557_out;
	wire [31:0] r558_out;
	wire [31:0] r559_out;
	wire [31:0] r560_out;
	wire [31:0] r561_out;
	wire [31:0] r562_out;
	wire [31:0] r563_out;
	wire [31:0] r564_out;
	wire [31:0] r565_out;
	wire [31:0] r566_out;
	wire [31:0] r567_out;
	wire [31:0] r568_out;
	wire [31:0] r569_out;
	wire [31:0] r570_out;
	wire [31:0] r571_out;
	wire [31:0] r572_out;
	wire [31:0] r573_out;
	wire [31:0] r574_out;
	wire [31:0] r575_out;
	wire [31:0] r576_out;
	wire [31:0] r577_out;
	wire [31:0] r578_out;
	wire [31:0] r579_out;
	wire [31:0] r580_out;
	wire [31:0] r581_out;
	wire [31:0] r582_out;
	wire [31:0] r583_out;
	wire [31:0] r584_out;
	wire [31:0] r585_out;
	wire [31:0] r586_out;
	wire [31:0] r587_out;
	wire [31:0] r588_out;
	wire [31:0] r589_out;
	wire [31:0] r590_out;
	wire [31:0] r591_out;
	wire [31:0] r592_out;
	wire [31:0] r593_out;
	wire [31:0] r594_out;
	wire [31:0] r595_out;
	wire [31:0] r596_out;
	wire [31:0] r597_out;
	wire [31:0] r598_out;
	wire [31:0] r599_out;
	wire [31:0] r600_out;
	wire [31:0] r601_out;
	wire [31:0] r602_out;
	wire [31:0] r603_out;
	wire [31:0] r604_out;
	wire [31:0] r605_out;
	wire [31:0] r606_out;
	wire [31:0] r607_out;
	wire [31:0] r608_out;
	wire [31:0] r609_out;
	wire [31:0] r610_out;
	wire [31:0] r611_out;
	wire [31:0] r612_out;
	wire [31:0] r613_out;
	wire [31:0] r614_out;
	wire [31:0] r615_out;
	wire [31:0] r616_out;
	wire [31:0] r617_out;
	wire [31:0] r618_out;
	wire [31:0] r619_out;
	wire [31:0] r620_out;
	wire [31:0] r621_out;
	wire [31:0] r622_out;
	wire [31:0] r623_out;
	wire [31:0] r624_out;
	wire [31:0] r625_out;
	wire [31:0] r626_out;
	wire [31:0] r627_out;
	wire [31:0] r628_out;
	wire [31:0] r629_out;
	wire [31:0] r630_out;
	wire [31:0] r631_out;
	wire [31:0] r632_out;
	wire [31:0] r633_out;
	wire [31:0] r634_out;
	wire [31:0] r635_out;
	wire [31:0] r636_out;
	wire [31:0] r637_out;
	wire [31:0] r638_out;
	wire [31:0] r639_out;
	wire [31:0] r640_out;
	wire [31:0] r641_out;
	wire [31:0] r642_out;
	wire [31:0] r643_out;
	wire [31:0] r644_out;
	wire [31:0] r645_out;
	wire [31:0] r646_out;
	wire [31:0] r647_out;
	wire [31:0] r648_out;
	wire [31:0] r649_out;
	wire [31:0] r650_out;
	wire [31:0] r651_out;
	wire [31:0] r652_out;
	wire [31:0] r653_out;
	wire [31:0] r654_out;
	wire [31:0] r655_out;
	wire [31:0] r656_out;
	wire [31:0] r657_out;
	wire [31:0] r658_out;
	wire [31:0] r659_out;
	wire [31:0] r660_out;
	wire [31:0] r661_out;
	wire [31:0] r662_out;
	wire [31:0] r663_out;
	wire [31:0] r664_out;
	wire [31:0] r665_out;
	wire [31:0] r666_out;
	wire [31:0] r667_out;
	wire [31:0] r668_out;
	wire [31:0] r669_out;
	wire [31:0] r670_out;
	wire [31:0] r671_out;
	wire [31:0] r672_out;
	wire [31:0] r673_out;
	wire [31:0] r674_out;
	wire [31:0] r675_out;
	wire [31:0] r676_out;
	wire [31:0] r677_out;
	wire [31:0] r678_out;
	wire [31:0] r679_out;
	wire [31:0] r680_out;
	wire [31:0] r681_out;
	wire [31:0] r682_out;
	wire [31:0] r683_out;
	wire [31:0] r684_out;
	wire [31:0] r685_out;
	wire [31:0] r686_out;
	wire [31:0] r687_out;
	wire [31:0] r688_out;
	wire [31:0] r689_out;
	wire [31:0] r690_out;
	wire [31:0] r691_out;
	wire [31:0] r692_out;
	wire [31:0] r693_out;
	wire [31:0] r694_out;
	wire [31:0] r695_out;
	wire [31:0] r696_out;
	wire [31:0] r697_out;
	wire [31:0] r698_out;
	wire [31:0] r699_out;
	wire [31:0] r700_out;
	wire [31:0] r701_out;
	wire [31:0] r702_out;
	wire [31:0] r703_out;
	wire [31:0] r704_out;
	wire [31:0] r705_out;
	wire [31:0] r706_out;
	wire [31:0] r707_out;
	wire [31:0] r708_out;
	wire [31:0] r709_out;
	wire [31:0] r710_out;
	wire [31:0] r711_out;
	wire [31:0] r712_out;
	wire [31:0] r713_out;
	wire [31:0] r714_out;
	wire [31:0] r715_out;
	wire [31:0] r716_out;
	wire [31:0] r717_out;
	wire [31:0] r718_out;
	wire [31:0] r719_out;
	wire [31:0] r720_out;
	wire [31:0] r721_out;
	wire [31:0] r722_out;
	wire [31:0] r723_out;
	wire [31:0] r724_out;
	wire [31:0] r725_out;
	wire [31:0] r726_out;
	wire [31:0] r727_out;
	wire [31:0] r728_out;
	wire [31:0] r729_out;
	wire [31:0] r730_out;
	wire [31:0] r731_out;
	wire [31:0] r732_out;
	wire [31:0] r733_out;
	wire [31:0] r734_out;
	wire [31:0] r735_out;
	wire [31:0] r736_out;
	wire [31:0] r737_out;
	wire [31:0] r738_out;
	wire [31:0] r739_out;
	wire [31:0] r740_out;
	wire [31:0] r741_out;
	wire [31:0] r742_out;
	wire [31:0] r743_out;
	wire [31:0] r744_out;
	wire [31:0] r745_out;
	wire [31:0] r746_out;
	wire [31:0] r747_out;
	wire [31:0] r748_out;
	wire [31:0] r749_out;
	wire [31:0] r750_out;
	wire [31:0] r751_out;
	wire [31:0] r752_out;
	wire [31:0] r753_out;
	wire [31:0] r754_out;
	wire [31:0] r755_out;
	wire [31:0] r756_out;
	wire [31:0] r757_out;
	wire [31:0] r758_out;
	wire [31:0] r759_out;
	wire [31:0] r760_out;
	wire [31:0] r761_out;
	wire [31:0] r762_out;
	wire [31:0] r763_out;
	wire [31:0] r764_out;
	wire [31:0] r765_out;
	wire [31:0] r766_out;
	wire [31:0] r767_out;
	wire [31:0] r768_out;
	wire [31:0] r769_out;
	wire [31:0] r770_out;
	wire [31:0] r771_out;
	wire [31:0] r772_out;
	wire [31:0] r773_out;
	wire [31:0] r774_out;
	wire [31:0] r775_out;
	wire [31:0] r776_out;
	wire [31:0] r777_out;
	wire [31:0] r778_out;
	wire [31:0] r779_out;
	wire [31:0] r780_out;
	wire [31:0] r781_out;
	wire [31:0] r782_out;
	wire [31:0] r783_out;
	wire [31:0] r784_out;
	wire [31:0] r785_out;
	wire [31:0] r786_out;
	wire [31:0] r787_out;
	wire [31:0] r788_out;
	wire [31:0] r789_out;
	wire [31:0] r790_out;
	wire [31:0] r791_out;
	wire [31:0] r792_out;
	wire [31:0] r793_out;
	wire [31:0] r794_out;
	wire [31:0] r795_out;
	wire [31:0] r796_out;
	wire [31:0] r797_out;
	wire [31:0] r798_out;
	wire [31:0] r799_out;
	wire [31:0] r800_out;
	wire [31:0] r801_out;
	wire [31:0] r802_out;
	wire [31:0] r803_out;
	wire [31:0] r804_out;
	wire [31:0] r805_out;
	wire [31:0] r806_out;
	wire [31:0] r807_out;
	wire [31:0] r808_out;
	wire [31:0] r809_out;
	wire [31:0] r810_out;
	wire [31:0] r811_out;
	wire [31:0] r812_out;
	wire [31:0] r813_out;
	wire [31:0] r814_out;
	wire [31:0] r815_out;
	wire [31:0] r816_out;
	wire [31:0] r817_out;
	wire [31:0] r818_out;
	wire [31:0] r819_out;
	wire [31:0] r820_out;
	wire [31:0] r821_out;
	wire [31:0] r822_out;
	wire [31:0] r823_out;
	wire [31:0] r824_out;
	wire [31:0] r825_out;
	wire [31:0] r826_out;
	wire [31:0] r827_out;
	wire [31:0] r828_out;
	wire [31:0] r829_out;
	wire [31:0] r830_out;
	wire [31:0] r831_out;
	wire [31:0] r832_out;
	wire [31:0] r833_out;
	wire [31:0] r834_out;
	wire [31:0] r835_out;
	wire [31:0] r836_out;
	wire [31:0] r837_out;
	wire [31:0] r838_out;
	wire [31:0] r839_out;
	wire [31:0] r840_out;
	wire [31:0] r841_out;
	wire [31:0] r842_out;
	wire [31:0] r843_out;
	wire [31:0] r844_out;
	wire [31:0] r845_out;
	wire [31:0] r846_out;
	wire [31:0] r847_out;
	wire [31:0] r848_out;
	wire [31:0] r849_out;
	wire [31:0] r850_out;
	wire [31:0] r851_out;
	wire [31:0] r852_out;
	wire [31:0] r853_out;
	wire [31:0] r854_out;
	wire [31:0] r855_out;
	wire [31:0] r856_out;
	wire [31:0] r857_out;
	wire [31:0] r858_out;
	wire [31:0] r859_out;
	wire [31:0] r860_out;
	wire [31:0] r861_out;
	wire [31:0] r862_out;
	wire [31:0] r863_out;
	wire [31:0] r864_out;
	wire [31:0] r865_out;
	wire [31:0] r866_out;
	wire [31:0] r867_out;
	wire [31:0] r868_out;
	wire [31:0] r869_out;
	wire [31:0] r870_out;
	wire [31:0] r871_out;
	wire [31:0] r872_out;
	wire [31:0] r873_out;
	wire [31:0] r874_out;
	wire [31:0] r875_out;
	wire [31:0] r876_out;
	wire [31:0] r877_out;
	wire [31:0] r878_out;
	wire [31:0] r879_out;
	wire [31:0] r880_out;
	wire [31:0] r881_out;
	wire [31:0] r882_out;
	wire [31:0] r883_out;
	wire [31:0] r884_out;
	wire [31:0] r885_out;
	wire [31:0] r886_out;
	wire [31:0] r887_out;
	wire [31:0] r888_out;
	wire [31:0] r889_out;
	wire [31:0] r890_out;
	wire [31:0] r891_out;
	wire [31:0] r892_out;
	wire [31:0] r893_out;
	wire [31:0] r894_out;
	wire [31:0] r895_out;
	wire [31:0] r896_out;
	wire [31:0] r897_out;
	wire [31:0] r898_out;
	wire [31:0] r899_out;
	wire [31:0] r900_out;
	wire [31:0] r901_out;
	wire [31:0] r902_out;
	wire [31:0] r903_out;
	wire [31:0] r904_out;
	wire [31:0] r905_out;
	wire [31:0] r906_out;
	wire [31:0] r907_out;
	wire [31:0] r908_out;
	wire [31:0] r909_out;
	wire [31:0] r910_out;
	wire [31:0] r911_out;
	wire [31:0] r912_out;
	wire [31:0] r913_out;
	wire [31:0] r914_out;
	wire [31:0] r915_out;
	wire [31:0] r916_out;
	wire [31:0] r917_out;
	wire [31:0] r918_out;
	wire [31:0] r919_out;
	wire [31:0] r920_out;
	wire [31:0] r921_out;
	wire [31:0] r922_out;
	wire [31:0] r923_out;
	wire [31:0] r924_out;
	wire [31:0] r925_out;
	wire [31:0] r926_out;
	wire [31:0] r927_out;
	wire [31:0] r928_out;
	wire [31:0] r929_out;
	wire [31:0] r930_out;
	wire [31:0] r931_out;
	wire [31:0] r932_out;
	wire [31:0] r933_out;
	wire [31:0] r934_out;
	wire [31:0] r935_out;
	wire [31:0] r936_out;
	wire [31:0] r937_out;
	wire [31:0] r938_out;
	wire [31:0] r939_out;
	wire [31:0] r940_out;
	wire [31:0] r941_out;
	wire [31:0] r942_out;
	wire [31:0] r943_out;
	wire [31:0] r944_out;
	wire [31:0] r945_out;
	wire [31:0] r946_out;
	wire [31:0] r947_out;
	wire [31:0] r948_out;
	wire [31:0] r949_out;
	wire [31:0] r950_out;
	wire [31:0] r951_out;
	wire [31:0] r952_out;
	wire [31:0] r953_out;
	wire [31:0] r954_out;
	wire [31:0] r955_out;
	wire [31:0] r956_out;
	wire [31:0] r957_out;
	wire [31:0] r958_out;
	wire [31:0] r959_out;
	wire [31:0] r960_out;
	wire [31:0] r961_out;
	wire [31:0] r962_out;
	wire [31:0] r963_out;
	wire [31:0] r964_out;
	wire [31:0] r965_out;
	wire [31:0] r966_out;
	wire [31:0] r967_out;
	wire [31:0] r968_out;
	wire [31:0] r969_out;
	wire [31:0] r970_out;
	wire [31:0] r971_out;
	wire [31:0] r972_out;
	wire [31:0] r973_out;
	wire [31:0] r974_out;
	wire [31:0] r975_out;
	wire [31:0] r976_out;
	wire [31:0] r977_out;
	wire [31:0] r978_out;
	wire [31:0] r979_out;
	wire [31:0] r980_out;
	wire [31:0] r981_out;
	wire [31:0] r982_out;
	wire [31:0] r983_out;
	wire [31:0] r984_out;
	wire [31:0] r985_out;
	wire [31:0] r986_out;
	wire [31:0] r987_out;
	wire [31:0] r988_out;
	wire [31:0] r989_out;
	wire [31:0] r990_out;
	wire [31:0] r991_out;
	wire [31:0] r992_out;
	wire [31:0] r993_out;
	wire [31:0] r994_out;
	wire [31:0] r995_out;
	wire [31:0] r996_out;
	wire [31:0] r997_out;
	wire [31:0] r998_out;
	wire [31:0] r999_out;
	wire [31:0] r1000_out;
	wire [31:0] r1001_out;
	wire [31:0] r1002_out;
	wire [31:0] r1003_out;
	wire [31:0] r1004_out;
	wire [31:0] r1005_out;
	wire [31:0] r1006_out;
	wire [31:0] r1007_out;
	wire [31:0] r1008_out;
	wire [31:0] r1009_out;
	wire [31:0] r1010_out;
	wire [31:0] r1011_out;
	wire [31:0] r1012_out;
	wire [31:0] r1013_out;
	wire [31:0] r1014_out;
	wire [31:0] r1015_out;
	wire [31:0] r1016_out;
	wire [31:0] r1017_out;
	wire [31:0] r1018_out;
	wire [31:0] r1019_out;
	wire [31:0] r1020_out;
	wire [31:0] r1021_out;
	wire [31:0] r1022_out;
	wire [31:0] r1023_out;
	wire [31:0] r1024_out;
	wire [31:0] r1025_out;
	wire [31:0] r1026_out;
	wire [31:0] r1027_out;
	wire [31:0] r1028_out;
	wire [31:0] r1029_out;
	wire [31:0] r1030_out;
	wire [31:0] r1031_out;
	wire [31:0] r1032_out;
	wire [31:0] r1033_out;
	wire [31:0] r1034_out;
	wire [31:0] r1035_out;
	wire [31:0] r1036_out;
	wire [31:0] r1037_out;
	wire [31:0] r1038_out;
	wire [31:0] r1039_out;
	wire [31:0] r1040_out;
	wire [31:0] r1041_out;
	wire [31:0] r1042_out;
	wire [31:0] r1043_out;
	wire [31:0] r1044_out;
	wire [31:0] r1045_out;
	wire [31:0] r1046_out;
	wire [31:0] r1047_out;
	wire [31:0] r1048_out;
	wire [31:0] r1049_out;
	wire [31:0] r1050_out;
	wire [31:0] r1051_out;
	wire [31:0] r1052_out;
	wire [31:0] r1053_out;
	wire [31:0] r1054_out;
	wire [31:0] r1055_out;
	wire [31:0] r1056_out;
	wire [31:0] r1057_out;
	wire [31:0] r1058_out;
	wire [31:0] r1059_out;
	wire [31:0] r1060_out;
	wire [31:0] r1061_out;
	wire [31:0] r1062_out;
	wire [31:0] r1063_out;
	wire [31:0] r1064_out;
	wire [31:0] r1065_out;
	wire [31:0] r1066_out;
	wire [31:0] r1067_out;
	wire [31:0] r1068_out;
	wire [31:0] r1069_out;
	wire [31:0] r1070_out;
	wire [31:0] r1071_out;
	wire [31:0] r1072_out;
	wire [31:0] r1073_out;
	wire [31:0] r1074_out;
	wire [31:0] r1075_out;
	wire [31:0] r1076_out;
	wire [31:0] r1077_out;
	wire [31:0] r1078_out;
	wire [31:0] r1079_out;
	wire [31:0] r1080_out;
	wire [31:0] r1081_out;
	wire [31:0] r1082_out;
	wire [31:0] r1083_out;
	wire [31:0] r1084_out;
	wire [31:0] r1085_out;
	wire [31:0] r1086_out;
	wire [31:0] r1087_out;
	wire [31:0] r1088_out;
	wire [31:0] r1089_out;
	wire [31:0] r1090_out;
	wire [31:0] r1091_out;
	wire [31:0] r1092_out;
	wire [31:0] r1093_out;
	wire [31:0] r1094_out;
	wire [31:0] r1095_out;
	wire [31:0] r1096_out;
	wire [31:0] r1097_out;
	wire [31:0] r1098_out;
	wire [31:0] r1099_out;
	wire [31:0] r1100_out;
	wire [31:0] r1101_out;
	wire [31:0] r1102_out;
	wire [31:0] r1103_out;
	wire [31:0] r1104_out;
	wire [31:0] r1105_out;
	wire [31:0] r1106_out;
	wire [31:0] r1107_out;
	wire [31:0] r1108_out;
	wire [31:0] r1109_out;
	wire [31:0] r1110_out;
	wire [31:0] r1111_out;
	wire [31:0] r1112_out;
	wire [31:0] r1113_out;
	wire [31:0] r1114_out;
	wire [31:0] r1115_out;
	wire [31:0] r1116_out;
	wire [31:0] r1117_out;
	wire [31:0] r1118_out;
	wire [31:0] r1119_out;
	wire [31:0] r1120_out;
	wire [31:0] r1121_out;
	wire [31:0] r1122_out;
	wire [31:0] r1123_out;
	wire [31:0] r1124_out;
	wire [31:0] r1125_out;
	wire [31:0] r1126_out;
	wire [31:0] r1127_out;
	wire [31:0] r1128_out;
	wire [31:0] r1129_out;
	wire [31:0] r1130_out;
	wire [31:0] r1131_out;
	wire [31:0] r1132_out;
	wire [31:0] r1133_out;
	wire [31:0] r1134_out;
	wire [31:0] r1135_out;
	wire [31:0] r1136_out;
	wire [31:0] r1137_out;
	wire [31:0] r1138_out;
	wire [31:0] r1139_out;
	wire [31:0] r1140_out;
	wire [31:0] r1141_out;
	wire [31:0] r1142_out;
	wire [31:0] r1143_out;
	wire [31:0] r1144_out;
	wire [31:0] r1145_out;
	wire [31:0] r1146_out;
	wire [31:0] r1147_out;
	wire [31:0] r1148_out;
	wire [31:0] r1149_out;
	wire [31:0] r1150_out;
	wire [31:0] r1151_out;
	wire [31:0] r1152_out;
	wire [31:0] r1153_out;
	wire [31:0] r1154_out;
	wire [31:0] r1155_out;
	wire [31:0] r1156_out;
	wire [31:0] r1157_out;
	wire [31:0] r1158_out;
	wire [31:0] r1159_out;
	wire [31:0] r1160_out;
	wire [31:0] r1161_out;
	wire [31:0] r1162_out;
	wire [31:0] r1163_out;
	wire [31:0] r1164_out;
	wire [31:0] r1165_out;
	wire [31:0] r1166_out;
	wire [31:0] r1167_out;
	wire [31:0] r1168_out;
	wire [31:0] r1169_out;
	wire [31:0] r1170_out;
	wire [31:0] r1171_out;
	wire [31:0] r1172_out;
	wire [31:0] r1173_out;
	wire [31:0] r1174_out;
	wire [31:0] r1175_out;
	wire [31:0] r1176_out;
	wire [31:0] r1177_out;
	wire [31:0] r1178_out;
	wire [31:0] r1179_out;
	wire [31:0] r1180_out;
	wire [31:0] r1181_out;
	wire [31:0] r1182_out;
	wire [31:0] r1183_out;
	wire [31:0] r1184_out;
	wire [31:0] r1185_out;
	wire [31:0] r1186_out;
	wire [31:0] r1187_out;
	wire [31:0] r1188_out;
	wire [31:0] r1189_out;
	wire [31:0] r1190_out;
	wire [31:0] r1191_out;
	wire [31:0] r1192_out;
	wire [31:0] r1193_out;
	wire [31:0] r1194_out;
	wire [31:0] r1195_out;
	wire [31:0] r1196_out;
	wire [31:0] r1197_out;
	wire [31:0] r1198_out;
	wire [31:0] r1199_out;
	wire [31:0] r1200_out;
	wire [31:0] r1201_out;
	wire [31:0] r1202_out;
	wire [31:0] r1203_out;
	wire [31:0] r1204_out;
	wire [31:0] r1205_out;
	wire [31:0] r1206_out;
	wire [31:0] r1207_out;
	wire [31:0] r1208_out;
	wire [31:0] r1209_out;
	wire [31:0] r1210_out;
	wire [31:0] r1211_out;
	wire [31:0] r1212_out;
	wire [31:0] r1213_out;
	wire [31:0] r1214_out;
	wire [31:0] r1215_out;
	wire [31:0] r1216_out;
	wire [31:0] r1217_out;
	wire [31:0] r1218_out;
	wire [31:0] r1219_out;
	wire [31:0] r1220_out;
	wire [31:0] r1221_out;
	wire [31:0] r1222_out;
	wire [31:0] r1223_out;
	wire [31:0] r1224_out;
	wire [31:0] r1225_out;
	wire [31:0] r1226_out;
	wire [31:0] r1227_out;
	wire [31:0] r1228_out;
	wire [31:0] r1229_out;
	wire [31:0] r1230_out;
	wire [31:0] r1231_out;
	wire [31:0] r1232_out;
	wire [31:0] r1233_out;
	wire [31:0] r1234_out;
	wire [31:0] r1235_out;
	wire [31:0] r1236_out;
	wire [31:0] r1237_out;
	wire [31:0] r1238_out;
	wire [31:0] r1239_out;
	wire [31:0] r1240_out;
	wire [31:0] r1241_out;
	wire [31:0] r1242_out;
	wire [31:0] r1243_out;
	wire [31:0] r1244_out;
	wire [31:0] r1245_out;
	wire [31:0] r1246_out;
	wire [31:0] r1247_out;
	wire [31:0] r1248_out;
	wire [31:0] r1249_out;
	wire [31:0] r1250_out;
	wire [31:0] r1251_out;
	wire [31:0] r1252_out;
	wire [31:0] r1253_out;
	wire [31:0] r1254_out;
	wire [31:0] r1255_out;
	wire [31:0] r1256_out;
	wire [31:0] r1257_out;
	wire [31:0] r1258_out;
	wire [31:0] r1259_out;
	wire [31:0] r1260_out;
	wire [31:0] r1261_out;
	wire [31:0] r1262_out;
	wire [31:0] r1263_out;
	wire [31:0] r1264_out;
	wire [31:0] r1265_out;
	wire [31:0] r1266_out;
	wire [31:0] r1267_out;
	wire [31:0] r1268_out;
	wire [31:0] r1269_out;
	wire [31:0] r1270_out;
	wire [31:0] r1271_out;
	wire [31:0] r1272_out;
	wire [31:0] r1273_out;
	wire [31:0] r1274_out;
	wire [31:0] r1275_out;
	wire [31:0] r1276_out;
	wire [31:0] r1277_out;
	wire [31:0] r1278_out;
	wire [31:0] r1279_out;
	wire [31:0] r1280_out;
	wire [31:0] r1281_out;
	wire [31:0] r1282_out;
	wire [31:0] r1283_out;
	wire [31:0] r1284_out;
	wire [31:0] r1285_out;
	wire [31:0] r1286_out;
	wire [31:0] r1287_out;
	wire [31:0] r1288_out;
	wire [31:0] r1289_out;
	wire [31:0] r1290_out;
	wire [31:0] r1291_out;
	wire [31:0] r1292_out;
	wire [31:0] r1293_out;
	wire [31:0] r1294_out;
	wire [31:0] r1295_out;
	wire [31:0] r1296_out;
	wire [31:0] r1297_out;
	wire [31:0] r1298_out;
	wire [31:0] r1299_out;
	wire [31:0] r1300_out;
	wire [31:0] r1301_out;
	wire [31:0] r1302_out;
	wire [31:0] r1303_out;
	wire [31:0] r1304_out;
	wire [31:0] r1305_out;
	wire [31:0] r1306_out;
	wire [31:0] r1307_out;
	wire [31:0] r1308_out;
	wire [31:0] r1309_out;
	wire [31:0] r1310_out;
	wire [31:0] r1311_out;
	wire [31:0] r1312_out;
	wire [31:0] r1313_out;
	wire [31:0] r1314_out;
	wire [31:0] r1315_out;
	wire [31:0] r1316_out;
	wire [31:0] r1317_out;
	wire [31:0] r1318_out;
	wire [31:0] r1319_out;
	wire [31:0] r1320_out;
	wire [31:0] r1321_out;
	wire [31:0] r1322_out;
	wire [31:0] r1323_out;
	wire [31:0] r1324_out;
	wire [31:0] r1325_out;
	wire [31:0] r1326_out;
	wire [31:0] r1327_out;
	wire [31:0] r1328_out;
	wire [31:0] r1329_out;
	wire [31:0] r1330_out;
	wire [31:0] r1331_out;
	wire [31:0] r1332_out;
	wire [31:0] r1333_out;
	wire [31:0] r1334_out;
	wire [31:0] r1335_out;
	wire [31:0] r1336_out;
	wire [31:0] r1337_out;
	wire [31:0] r1338_out;
	wire [31:0] r1339_out;
	wire [31:0] r1340_out;
	wire [31:0] r1341_out;
	wire [31:0] r1342_out;
	wire [31:0] r1343_out;
	wire [31:0] r1344_out;
	wire [31:0] r1345_out;
	wire [31:0] r1346_out;
	wire [31:0] r1347_out;
	wire [31:0] r1348_out;
	wire [31:0] r1349_out;
	wire [31:0] r1350_out;
	wire [31:0] r1351_out;
	wire [31:0] r1352_out;
	wire [31:0] r1353_out;
	wire [31:0] r1354_out;
	wire [31:0] r1355_out;
	wire [31:0] r1356_out;
	wire [31:0] r1357_out;
	wire [31:0] r1358_out;
	wire [31:0] r1359_out;
	wire [31:0] r1360_out;
	wire [31:0] r1361_out;
	wire [31:0] r1362_out;
	wire [31:0] r1363_out;
	wire [31:0] r1364_out;
	wire [31:0] r1365_out;
	wire [31:0] r1366_out;
	wire [31:0] r1367_out;
	wire [31:0] r1368_out;
	wire [31:0] r1369_out;
	wire [31:0] r1370_out;
	wire [31:0] r1371_out;
	wire [31:0] r1372_out;
	wire [31:0] r1373_out;
	wire [31:0] r1374_out;
	wire [31:0] r1375_out;
	wire [31:0] r1376_out;
	wire [31:0] r1377_out;
	wire [31:0] r1378_out;
	wire [31:0] r1379_out;
	wire [31:0] r1380_out;
	wire [31:0] r1381_out;
	wire [31:0] r1382_out;
	wire [31:0] r1383_out;
	wire [31:0] r1384_out;
	wire [31:0] r1385_out;
	wire [31:0] r1386_out;
	wire [31:0] r1387_out;
	wire [31:0] r1388_out;
	wire [31:0] r1389_out;
	wire [31:0] r1390_out;
	wire [31:0] r1391_out;
	wire [31:0] r1392_out;
	wire [31:0] r1393_out;
	wire [31:0] r1394_out;
	wire [31:0] r1395_out;
	wire [31:0] r1396_out;
	wire [31:0] r1397_out;
	wire [31:0] r1398_out;
	wire [31:0] r1399_out;
	wire [31:0] r1400_out;
	wire [31:0] r1401_out;
	wire [31:0] r1402_out;
	wire [31:0] r1403_out;
	wire [31:0] r1404_out;
	wire [31:0] r1405_out;
	wire [31:0] r1406_out;
	wire [31:0] r1407_out;
	wire [31:0] r1408_out;
	wire [31:0] r1409_out;
	wire [31:0] r1410_out;
	wire [31:0] r1411_out;
	wire [31:0] r1412_out;
	wire [31:0] r1413_out;
	wire [31:0] r1414_out;
	wire [31:0] r1415_out;
	wire [31:0] r1416_out;
	wire [31:0] r1417_out;
	wire [31:0] r1418_out;
	wire [31:0] r1419_out;
	wire [31:0] r1420_out;
	wire [31:0] r1421_out;
	wire [31:0] r1422_out;
	wire [31:0] r1423_out;
	wire [31:0] r1424_out;
	wire [31:0] r1425_out;
	wire [31:0] r1426_out;
	wire [31:0] r1427_out;
	wire [31:0] r1428_out;
	wire [31:0] r1429_out;
	wire [31:0] r1430_out;
	wire [31:0] r1431_out;
	wire [31:0] r1432_out;
	wire [31:0] r1433_out;
	wire [31:0] r1434_out;
	wire [31:0] r1435_out;
	wire [31:0] r1436_out;
	wire [31:0] r1437_out;
	wire [31:0] r1438_out;
	wire [31:0] r1439_out;
	wire [31:0] r1440_out;
	wire [31:0] r1441_out;
	wire [31:0] r1442_out;
	wire [31:0] r1443_out;
	wire [31:0] r1444_out;
	wire [31:0] r1445_out;
	wire [31:0] r1446_out;
	wire [31:0] r1447_out;
	wire [31:0] r1448_out;
	wire [31:0] r1449_out;
	wire [31:0] r1450_out;
	wire [31:0] r1451_out;
	wire [31:0] r1452_out;
	wire [31:0] r1453_out;
	wire [31:0] r1454_out;
	wire [31:0] r1455_out;
	wire [31:0] r1456_out;
	wire [31:0] r1457_out;
	wire [31:0] r1458_out;
	wire [31:0] r1459_out;
	wire [31:0] r1460_out;
	wire [31:0] r1461_out;
	wire [31:0] r1462_out;
	wire [31:0] r1463_out;
	wire [31:0] r1464_out;
	wire [31:0] r1465_out;
	wire [31:0] r1466_out;
	wire [31:0] r1467_out;
	wire [31:0] r1468_out;
	wire [31:0] r1469_out;
	wire [31:0] r1470_out;
	wire [31:0] r1471_out;
	wire [31:0] r1472_out;
	wire [31:0] r1473_out;
	wire [31:0] r1474_out;
	wire [31:0] r1475_out;
	wire [31:0] r1476_out;
	wire [31:0] r1477_out;
	wire [31:0] r1478_out;
	wire [31:0] r1479_out;
	wire [31:0] r1480_out;
	wire [31:0] r1481_out;
	wire [31:0] r1482_out;
	wire [31:0] r1483_out;
	wire [31:0] r1484_out;
	wire [31:0] r1485_out;
	wire [31:0] r1486_out;
	wire [31:0] r1487_out;
	wire [31:0] r1488_out;
	wire [31:0] r1489_out;
	wire [31:0] r1490_out;
	wire [31:0] r1491_out;
	wire [31:0] r1492_out;
	wire [31:0] r1493_out;
	wire [31:0] r1494_out;
	wire [31:0] r1495_out;
	wire [31:0] r1496_out;
	wire [31:0] r1497_out;
	wire [31:0] r1498_out;
	wire [31:0] r1499_out;
	wire [31:0] r1500_out;
	wire [31:0] r1501_out;
	wire [31:0] r1502_out;
	wire [31:0] r1503_out;
	wire [31:0] r1504_out;
	wire [31:0] r1505_out;
	wire [31:0] r1506_out;
	wire [31:0] r1507_out;
	wire [31:0] r1508_out;
	wire [31:0] r1509_out;
	wire [31:0] r1510_out;
	wire [31:0] r1511_out;
	wire [31:0] r1512_out;
	wire [31:0] r1513_out;
	wire [31:0] r1514_out;
	wire [31:0] r1515_out;
	wire [31:0] r1516_out;
	wire [31:0] r1517_out;
	wire [31:0] r1518_out;
	wire [31:0] r1519_out;
	wire [31:0] r1520_out;
	wire [31:0] r1521_out;
	wire [31:0] r1522_out;
	wire [31:0] r1523_out;
	wire [31:0] r1524_out;
	wire [31:0] r1525_out;
	wire [31:0] r1526_out;
	wire [31:0] r1527_out;
	wire [31:0] r1528_out;
	wire [31:0] r1529_out;
	wire [31:0] r1530_out;
	wire [31:0] r1531_out;
	wire [31:0] r1532_out;
	wire [31:0] r1533_out;
	wire [31:0] r1534_out;
	wire [31:0] r1535_out;
	wire [31:0] r1536_out;
	wire [31:0] r1537_out;
	wire [31:0] r1538_out;
	wire [31:0] r1539_out;
	wire [31:0] r1540_out;
	wire [31:0] r1541_out;
	wire [31:0] r1542_out;
	wire [31:0] r1543_out;
	wire [31:0] r1544_out;
	wire [31:0] r1545_out;
	wire [31:0] r1546_out;
	wire [31:0] r1547_out;
	wire [31:0] r1548_out;
	wire [31:0] r1549_out;
	wire [31:0] r1550_out;
	wire [31:0] r1551_out;
	wire [31:0] r1552_out;
	wire [31:0] r1553_out;
	wire [31:0] r1554_out;
	wire [31:0] r1555_out;
	wire [31:0] r1556_out;
	wire [31:0] r1557_out;
	wire [31:0] r1558_out;
	wire [31:0] r1559_out;
	wire [31:0] r1560_out;
	wire [31:0] r1561_out;
	wire [31:0] r1562_out;
	wire [31:0] r1563_out;
	wire [31:0] r1564_out;
	wire [31:0] r1565_out;
	wire [31:0] r1566_out;
	wire [31:0] r1567_out;
	wire [31:0] r1568_out;
	wire [31:0] r1569_out;
	wire [31:0] r1570_out;
	wire [31:0] r1571_out;
	wire [31:0] r1572_out;
	wire [31:0] r1573_out;
	wire [31:0] r1574_out;
	wire [31:0] r1575_out;
	wire [31:0] r1576_out;
	wire [31:0] r1577_out;
	wire [31:0] r1578_out;
	wire [31:0] r1579_out;
	wire [31:0] r1580_out;
	wire [31:0] r1581_out;
	wire [31:0] r1582_out;
	wire [31:0] r1583_out;
	wire [31:0] r1584_out;
	wire [31:0] r1585_out;
	wire [31:0] r1586_out;
	wire [31:0] r1587_out;
	wire [31:0] r1588_out;
	wire [31:0] r1589_out;
	wire [31:0] r1590_out;
	wire [31:0] r1591_out;
	wire [31:0] r1592_out;
	wire [31:0] r1593_out;
	wire [31:0] r1594_out;
	wire [31:0] r1595_out;
	wire [31:0] r1596_out;
	wire [31:0] r1597_out;
	wire [31:0] r1598_out;
	wire [31:0] r1599_out;
	wire [31:0] r1600_out;
	wire [31:0] r1601_out;
	wire [31:0] r1602_out;
	wire [31:0] r1603_out;
	wire [31:0] r1604_out;
	wire [31:0] r1605_out;
	wire [31:0] r1606_out;
	wire [31:0] r1607_out;
	wire [31:0] r1608_out;
	wire [31:0] r1609_out;
	wire [31:0] r1610_out;
	wire [31:0] r1611_out;
	wire [31:0] r1612_out;
	wire [31:0] r1613_out;
	wire [31:0] r1614_out;
	wire [31:0] r1615_out;
	wire [31:0] r1616_out;
	wire [31:0] r1617_out;
	wire [31:0] r1618_out;
	wire [31:0] r1619_out;
	wire [31:0] r1620_out;
	wire [31:0] r1621_out;
	wire [31:0] r1622_out;
	wire [31:0] r1623_out;
	wire [31:0] r1624_out;
	wire [31:0] r1625_out;
	wire [31:0] r1626_out;
	wire [31:0] r1627_out;
	wire [31:0] r1628_out;
	wire [31:0] r1629_out;
	wire [31:0] r1630_out;
	wire [31:0] r1631_out;
	wire [31:0] r1632_out;
	wire [31:0] r1633_out;
	wire [31:0] r1634_out;
	wire [31:0] r1635_out;
	wire [31:0] r1636_out;
	wire [31:0] r1637_out;
	wire [31:0] r1638_out;
	wire [31:0] r1639_out;
	wire [31:0] r1640_out;
	wire [31:0] r1641_out;
	wire [31:0] r1642_out;
	wire [31:0] r1643_out;
	wire [31:0] r1644_out;
	wire [31:0] r1645_out;
	wire [31:0] r1646_out;
	wire [31:0] r1647_out;
	wire [31:0] r1648_out;
	wire [31:0] r1649_out;
	wire [31:0] r1650_out;
	wire [31:0] r1651_out;
	wire [31:0] r1652_out;
	wire [31:0] r1653_out;
	wire [31:0] r1654_out;
	wire [31:0] r1655_out;
	wire [31:0] r1656_out;
	wire [31:0] r1657_out;
	wire [31:0] r1658_out;
	wire [31:0] r1659_out;
	wire [31:0] r1660_out;
	wire [31:0] r1661_out;
	wire [31:0] r1662_out;
	wire [31:0] r1663_out;
	wire [31:0] r1664_out;
	wire [31:0] r1665_out;
	wire [31:0] r1666_out;
	wire [31:0] r1667_out;
	wire [31:0] r1668_out;
	wire [31:0] r1669_out;
	wire [31:0] r1670_out;
	wire [31:0] r1671_out;
	wire [31:0] r1672_out;
	wire [31:0] r1673_out;
	wire [31:0] r1674_out;
	wire [31:0] r1675_out;
	wire [31:0] r1676_out;
	wire [31:0] r1677_out;
	wire [31:0] r1678_out;
	wire [31:0] r1679_out;
	wire [31:0] r1680_out;
	wire [31:0] r1681_out;
	wire [31:0] r1682_out;
	wire [31:0] r1683_out;
	wire [31:0] r1684_out;
	wire [31:0] r1685_out;
	wire [31:0] r1686_out;
	wire [31:0] r1687_out;
	wire [31:0] r1688_out;
	wire [31:0] r1689_out;
	wire [31:0] r1690_out;
	wire [31:0] r1691_out;
	wire [31:0] r1692_out;
	wire [31:0] r1693_out;
	wire [31:0] r1694_out;
	wire [31:0] r1695_out;
	wire [31:0] r1696_out;
	wire [31:0] r1697_out;
	wire [31:0] r1698_out;
	wire [31:0] r1699_out;
	wire [31:0] r1700_out;
	wire [31:0] r1701_out;
	wire [31:0] r1702_out;
	wire [31:0] r1703_out;
	wire [31:0] r1704_out;
	wire [31:0] r1705_out;
	wire [31:0] r1706_out;
	wire [31:0] r1707_out;
	wire [31:0] r1708_out;
	wire [31:0] r1709_out;
	wire [31:0] r1710_out;
	wire [31:0] r1711_out;
	wire [31:0] r1712_out;
	wire [31:0] r1713_out;
	wire [31:0] r1714_out;
	wire [31:0] r1715_out;
	wire [31:0] r1716_out;
	wire [31:0] r1717_out;
	wire [31:0] r1718_out;
	wire [31:0] r1719_out;
	wire [31:0] r1720_out;
	wire [31:0] r1721_out;
	wire [31:0] r1722_out;
	wire [31:0] r1723_out;
	wire [31:0] r1724_out;
	wire [31:0] r1725_out;
	wire [31:0] r1726_out;
	wire [31:0] r1727_out;
	wire [31:0] r1728_out;
	wire [31:0] r1729_out;
	wire [31:0] r1730_out;
	wire [31:0] r1731_out;
	wire [31:0] r1732_out;
	wire [31:0] r1733_out;
	wire [31:0] r1734_out;
	wire [31:0] r1735_out;
	wire [31:0] r1736_out;
	wire [31:0] r1737_out;
	wire [31:0] r1738_out;
	wire [31:0] r1739_out;
	wire [31:0] r1740_out;
	wire [31:0] r1741_out;
	wire [31:0] r1742_out;
	wire [31:0] r1743_out;
	wire [31:0] r1744_out;
	wire [31:0] r1745_out;
	wire [31:0] r1746_out;
	wire [31:0] r1747_out;
	wire [31:0] r1748_out;
	wire [31:0] r1749_out;
	wire [31:0] r1750_out;
	wire [31:0] r1751_out;
	wire [31:0] r1752_out;
	wire [31:0] r1753_out;
	wire [31:0] r1754_out;
	wire [31:0] r1755_out;
	wire [31:0] r1756_out;
	wire [31:0] r1757_out;
	wire [31:0] r1758_out;
	wire [31:0] r1759_out;
	wire [31:0] r1760_out;
	wire [31:0] r1761_out;
	wire [31:0] r1762_out;
	wire [31:0] r1763_out;
	wire [31:0] r1764_out;
	wire [31:0] r1765_out;
	wire [31:0] r1766_out;
	wire [31:0] r1767_out;
	wire [31:0] r1768_out;
	wire [31:0] r1769_out;
	wire [31:0] r1770_out;
	wire [31:0] r1771_out;
	wire [31:0] r1772_out;
	wire [31:0] r1773_out;
	wire [31:0] r1774_out;
	wire [31:0] r1775_out;
	wire [31:0] r1776_out;
	wire [31:0] r1777_out;
	wire [31:0] r1778_out;
	wire [31:0] r1779_out;
	wire [31:0] r1780_out;
	wire [31:0] r1781_out;
	wire [31:0] r1782_out;
	wire [31:0] r1783_out;
	wire [31:0] r1784_out;
	wire [31:0] r1785_out;
	wire [31:0] r1786_out;
	wire [31:0] r1787_out;
	wire [31:0] r1788_out;
	wire [31:0] r1789_out;
	wire [31:0] r1790_out;
	wire [31:0] r1791_out;
	wire [31:0] r1792_out;
	wire [31:0] r1793_out;
	wire [31:0] r1794_out;
	wire [31:0] r1795_out;
	wire [31:0] r1796_out;
	wire [31:0] r1797_out;
	wire [31:0] r1798_out;
	wire [31:0] r1799_out;
	wire [31:0] r1800_out;
	wire [31:0] r1801_out;
	wire [31:0] r1802_out;
	wire [31:0] r1803_out;
	wire [31:0] r1804_out;
	wire [31:0] r1805_out;
	wire [31:0] r1806_out;
	wire [31:0] r1807_out;
	wire [31:0] r1808_out;
	wire [31:0] r1809_out;
	wire [31:0] r1810_out;
	wire [31:0] r1811_out;
	wire [31:0] r1812_out;
	wire [31:0] r1813_out;
	wire [31:0] r1814_out;
	wire [31:0] r1815_out;
	wire [31:0] r1816_out;
	wire [31:0] r1817_out;
	wire [31:0] r1818_out;
	wire [31:0] r1819_out;
	wire [31:0] r1820_out;
	wire [31:0] r1821_out;
	wire [31:0] r1822_out;
	wire [31:0] r1823_out;
	wire [31:0] r1824_out;
	wire [31:0] r1825_out;
	wire [31:0] r1826_out;
	wire [31:0] r1827_out;
	wire [31:0] r1828_out;
	wire [31:0] r1829_out;
	wire [31:0] r1830_out;
	wire [31:0] r1831_out;
	wire [31:0] r1832_out;
	wire [31:0] r1833_out;
	wire [31:0] r1834_out;
	wire [31:0] r1835_out;
	wire [31:0] r1836_out;
	wire [31:0] r1837_out;
	wire [31:0] r1838_out;
	wire [31:0] r1839_out;
	wire [31:0] r1840_out;
	wire [31:0] r1841_out;
	wire [31:0] r1842_out;
	wire [31:0] r1843_out;
	wire [31:0] r1844_out;
	wire [31:0] r1845_out;
	wire [31:0] r1846_out;
	wire [31:0] r1847_out;
	wire [31:0] r1848_out;
	wire [31:0] r1849_out;
	wire [31:0] r1850_out;
	wire [31:0] r1851_out;
	wire [31:0] r1852_out;
	wire [31:0] r1853_out;
	wire [31:0] r1854_out;
	wire [31:0] r1855_out;
	wire [31:0] r1856_out;
	wire [31:0] r1857_out;
	wire [31:0] r1858_out;
	wire [31:0] r1859_out;
	wire [31:0] r1860_out;
	wire [31:0] r1861_out;
	wire [31:0] r1862_out;
	wire [31:0] r1863_out;
	wire [31:0] r1864_out;
	wire [31:0] r1865_out;
	wire [31:0] r1866_out;
	wire [31:0] r1867_out;
	wire [31:0] r1868_out;
	wire [31:0] r1869_out;
	wire [31:0] r1870_out;
	wire [31:0] r1871_out;
	wire [31:0] r1872_out;
	wire [31:0] r1873_out;
	wire [31:0] r1874_out;
	wire [31:0] r1875_out;
	wire [31:0] r1876_out;
	wire [31:0] r1877_out;
	wire [31:0] r1878_out;
	wire [31:0] r1879_out;
	wire [31:0] r1880_out;
	wire [31:0] r1881_out;
	wire [31:0] r1882_out;
	wire [31:0] r1883_out;
	wire [31:0] r1884_out;
	wire [31:0] r1885_out;
	wire [31:0] r1886_out;
	wire [31:0] r1887_out;
	wire [31:0] r1888_out;
	wire [31:0] r1889_out;
	wire [31:0] r1890_out;
	wire [31:0] r1891_out;
	wire [31:0] r1892_out;
	wire [31:0] r1893_out;
	wire [31:0] r1894_out;
	wire [31:0] r1895_out;
	wire [31:0] r1896_out;
	wire [31:0] r1897_out;
	wire [31:0] r1898_out;
	wire [31:0] r1899_out;
	wire [31:0] r1900_out;
	wire [31:0] r1901_out;
	wire [31:0] r1902_out;
	wire [31:0] r1903_out;
	wire [31:0] r1904_out;
	wire [31:0] r1905_out;
	wire [31:0] r1906_out;
	wire [31:0] r1907_out;
	wire [31:0] r1908_out;
	wire [31:0] r1909_out;
	wire [31:0] r1910_out;
	wire [31:0] r1911_out;
	wire [31:0] r1912_out;
	wire [31:0] r1913_out;
	wire [31:0] r1914_out;
	wire [31:0] r1915_out;
	wire [31:0] r1916_out;
	wire [31:0] r1917_out;
	wire [31:0] r1918_out;
	wire [31:0] r1919_out;
	wire [31:0] r1920_out;
	wire [31:0] r1921_out;
	wire [31:0] r1922_out;
	wire [31:0] r1923_out;
	wire [31:0] r1924_out;
	wire [31:0] r1925_out;
	wire [31:0] r1926_out;
	wire [31:0] r1927_out;
	wire [31:0] r1928_out;
	wire [31:0] r1929_out;
	wire [31:0] r1930_out;
	wire [31:0] r1931_out;
	wire [31:0] r1932_out;
	wire [31:0] r1933_out;
	wire [31:0] r1934_out;
	wire [31:0] r1935_out;
	wire [31:0] r1936_out;
	wire [31:0] r1937_out;
	wire [31:0] r1938_out;
	wire [31:0] r1939_out;
	wire [31:0] r1940_out;
	wire [31:0] r1941_out;
	wire [31:0] r1942_out;
	wire [31:0] r1943_out;
	wire [31:0] r1944_out;
	wire [31:0] r1945_out;
	wire [31:0] r1946_out;
	wire [31:0] r1947_out;
	wire [31:0] r1948_out;
	wire [31:0] r1949_out;
	wire [31:0] r1950_out;
	wire [31:0] r1951_out;
	wire [31:0] r1952_out;
	wire [31:0] r1953_out;
	wire [31:0] r1954_out;
	wire [31:0] r1955_out;
	wire [31:0] r1956_out;
	wire [31:0] r1957_out;
	wire [31:0] r1958_out;
	wire [31:0] r1959_out;
	wire [31:0] r1960_out;
	wire [31:0] r1961_out;
	wire [31:0] r1962_out;
	wire [31:0] r1963_out;
	wire [31:0] r1964_out;
	wire [31:0] r1965_out;
	wire [31:0] r1966_out;
	wire [31:0] r1967_out;
	wire [31:0] r1968_out;
	wire [31:0] r1969_out;
	wire [31:0] r1970_out;
	wire [31:0] r1971_out;
	wire [31:0] r1972_out;
	wire [31:0] r1973_out;
	wire [31:0] r1974_out;
	wire [31:0] r1975_out;
	wire [31:0] r1976_out;
	wire [31:0] r1977_out;
	wire [31:0] r1978_out;
	wire [31:0] r1979_out;
	wire [31:0] r1980_out;
	wire [31:0] r1981_out;
	wire [31:0] r1982_out;
	wire [31:0] r1983_out;
	wire [31:0] r1984_out;
	wire [31:0] r1985_out;
	wire [31:0] r1986_out;
	wire [31:0] r1987_out;
	wire [31:0] r1988_out;
	wire [31:0] r1989_out;
	wire [31:0] r1990_out;
	wire [31:0] r1991_out;
	wire [31:0] r1992_out;
	wire [31:0] r1993_out;
	wire [31:0] r1994_out;
	wire [31:0] r1995_out;
	wire [31:0] r1996_out;
	wire [31:0] r1997_out;
	wire [31:0] r1998_out;
	wire [31:0] r1999_out;
	wire [31:0] r2000_out;
	wire [31:0] r2001_out;
	wire [31:0] r2002_out;
	wire [31:0] r2003_out;
	wire [31:0] r2004_out;
	wire [31:0] r2005_out;
	wire [31:0] r2006_out;
	wire [31:0] r2007_out;
	wire [31:0] r2008_out;
	wire [31:0] r2009_out;
	wire [31:0] r2010_out;
	wire [31:0] r2011_out;
	wire [31:0] r2012_out;
	wire [31:0] r2013_out;
	wire [31:0] r2014_out;
	wire [31:0] r2015_out;
	wire [31:0] r2016_out;
	wire [31:0] r2017_out;
	wire [31:0] r2018_out;
	wire [31:0] r2019_out;
	wire [31:0] r2020_out;
	wire [31:0] r2021_out;
	wire [31:0] r2022_out;
	wire [31:0] r2023_out;
	wire [31:0] r2024_out;
	wire [31:0] r2025_out;
	wire [31:0] r2026_out;
	wire [31:0] r2027_out;
	wire [31:0] r2028_out;
	wire [31:0] r2029_out;
	wire [31:0] r2030_out;
	wire [31:0] r2031_out;
	wire [31:0] r2032_out;
	wire [31:0] r2033_out;
	wire [31:0] r2034_out;
	wire [31:0] r2035_out;
	wire [31:0] r2036_out;
	wire [31:0] r2037_out;
	wire [31:0] r2038_out;
	wire [31:0] r2039_out;
	wire [31:0] r2040_out;
	wire [31:0] r2041_out;
	wire [31:0] r2042_out;
	wire [31:0] r2043_out;
	wire [31:0] r2044_out;
	wire [31:0] r2045_out;
	wire [31:0] r2046_out;
	wire [31:0] r2047_out;
	wire [31:0] r2048_out;
	wire [31:0] r2049_out;
	wire [31:0] r2050_out;
	wire [31:0] r2051_out;
	wire [31:0] r2052_out;
	wire [31:0] r2053_out;
	wire [31:0] r2054_out;
	wire [31:0] r2055_out;
	wire [31:0] r2056_out;
	wire [31:0] r2057_out;
	wire [31:0] r2058_out;
	wire [31:0] r2059_out;
	wire [31:0] r2060_out;
	wire [31:0] r2061_out;
	wire [31:0] r2062_out;
	wire [31:0] r2063_out;
	wire [31:0] r2064_out;
	wire [31:0] r2065_out;
	wire [31:0] r2066_out;
	wire [31:0] r2067_out;
	wire [31:0] r2068_out;
	wire [31:0] r2069_out;
	wire [31:0] r2070_out;
	wire [31:0] r2071_out;
	wire [31:0] r2072_out;
	wire [31:0] r2073_out;
	wire [31:0] r2074_out;
	wire [31:0] r2075_out;
	wire [31:0] r2076_out;
	wire [31:0] r2077_out;
	wire [31:0] r2078_out;
	wire [31:0] r2079_out;
	wire [31:0] r2080_out;
	wire [31:0] r2081_out;
	wire [31:0] r2082_out;
	wire [31:0] r2083_out;
	wire [31:0] r2084_out;
	wire [31:0] r2085_out;
	wire [31:0] r2086_out;
	wire [31:0] r2087_out;
	wire [31:0] r2088_out;
	wire [31:0] r2089_out;
	wire [31:0] r2090_out;
	wire [31:0] r2091_out;
	wire [31:0] r2092_out;
	wire [31:0] r2093_out;
	wire [31:0] r2094_out;
	wire [31:0] r2095_out;
	wire [31:0] r2096_out;
	wire [31:0] r2097_out;
	wire [31:0] r2098_out;
	wire [31:0] r2099_out;
	wire [31:0] r2100_out;
	wire [31:0] r2101_out;
	wire [31:0] r2102_out;
	wire [31:0] r2103_out;
	wire [31:0] r2104_out;
	wire [31:0] r2105_out;
	wire [31:0] r2106_out;
	wire [31:0] r2107_out;
	wire [31:0] r2108_out;
	wire [31:0] r2109_out;
	wire [31:0] r2110_out;
	wire [31:0] r2111_out;
	wire [31:0] r2112_out;
	wire [31:0] r2113_out;
	wire [31:0] r2114_out;
	wire [31:0] r2115_out;
	wire [31:0] r2116_out;
	wire [31:0] r2117_out;
	wire [31:0] r2118_out;
	wire [31:0] r2119_out;
	wire [31:0] r2120_out;
	wire [31:0] r2121_out;
	wire [31:0] r2122_out;
	wire [31:0] r2123_out;
	wire [31:0] r2124_out;
	wire [31:0] r2125_out;
	wire [31:0] r2126_out;
	wire [31:0] r2127_out;
	wire [31:0] r2128_out;
	wire [31:0] r2129_out;
	wire [31:0] r2130_out;
	wire [31:0] r2131_out;
	wire [31:0] r2132_out;
	wire [31:0] r2133_out;
	wire [31:0] r2134_out;
	wire [31:0] r2135_out;
	wire [31:0] r2136_out;
	wire [31:0] r2137_out;
	wire [31:0] r2138_out;
	wire [31:0] r2139_out;
	wire [31:0] r2140_out;
	wire [31:0] r2141_out;
	wire [31:0] r2142_out;
	wire [31:0] r2143_out;
	wire [31:0] r2144_out;
	wire [31:0] r2145_out;
	wire [31:0] r2146_out;
	wire [31:0] r2147_out;
	wire [31:0] r2148_out;
	wire [31:0] r2149_out;
	wire [31:0] r2150_out;
	wire [31:0] r2151_out;
	wire [31:0] r2152_out;
	wire [31:0] r2153_out;
	wire [31:0] r2154_out;
	wire [31:0] r2155_out;
	wire [31:0] r2156_out;
	wire [31:0] r2157_out;
	wire [31:0] r2158_out;
	wire [31:0] r2159_out;
	wire [31:0] r2160_out;
	wire [31:0] r2161_out;
	wire [31:0] r2162_out;
	wire [31:0] r2163_out;
	wire [31:0] r2164_out;
	wire [31:0] r2165_out;
	wire [31:0] r2166_out;
	wire [31:0] r2167_out;
	wire [31:0] r2168_out;
	wire [31:0] r2169_out;
	wire [31:0] r2170_out;
	wire [31:0] r2171_out;
	wire [31:0] r2172_out;
	wire [31:0] r2173_out;
	wire [31:0] r2174_out;
	wire [31:0] r2175_out;
	wire [31:0] r2176_out;
	wire [31:0] r2177_out;
	wire [31:0] r2178_out;
	wire [31:0] r2179_out;
	wire [31:0] r2180_out;
	wire [31:0] r2181_out;
	wire [31:0] r2182_out;
	wire [31:0] r2183_out;
	wire [31:0] r2184_out;
	wire [31:0] r2185_out;
	wire [31:0] r2186_out;
	wire [31:0] r2187_out;
	wire [31:0] r2188_out;
	wire [31:0] r2189_out;
	wire [31:0] r2190_out;
	wire [31:0] r2191_out;
	wire [31:0] r2192_out;
	wire [31:0] r2193_out;
	wire [31:0] r2194_out;
	wire [31:0] r2195_out;
	wire [31:0] r2196_out;
	wire [31:0] r2197_out;
	wire [31:0] r2198_out;
	wire [31:0] r2199_out;
	wire [31:0] r2200_out;
	wire [31:0] r2201_out;
	wire [31:0] r2202_out;
	wire [31:0] r2203_out;
	wire [31:0] r2204_out;
	wire [31:0] r2205_out;
	wire [31:0] r2206_out;
	wire [31:0] r2207_out;
	wire [31:0] r2208_out;
	wire [31:0] r2209_out;
	wire [31:0] r2210_out;
	wire [31:0] r2211_out;
	wire [31:0] r2212_out;
	wire [31:0] r2213_out;
	wire [31:0] r2214_out;
	wire [31:0] r2215_out;
	wire [31:0] r2216_out;
	wire [31:0] r2217_out;
	wire [31:0] r2218_out;
	wire [31:0] r2219_out;
	wire [31:0] r2220_out;
	wire [31:0] r2221_out;
	wire [31:0] r2222_out;
	wire [31:0] r2223_out;
	wire [31:0] r2224_out;
	wire [31:0] r2225_out;
	wire [31:0] r2226_out;
	wire [31:0] r2227_out;
	wire [31:0] r2228_out;
	wire [31:0] r2229_out;
	wire [31:0] r2230_out;
	wire [31:0] r2231_out;
	wire [31:0] r2232_out;
	wire [31:0] r2233_out;
	wire [31:0] r2234_out;
	wire [31:0] r2235_out;
	wire [31:0] r2236_out;
	wire [31:0] r2237_out;
	wire [31:0] r2238_out;
	wire [31:0] r2239_out;
	wire [31:0] r2240_out;
	wire [31:0] r2241_out;
	wire [31:0] r2242_out;
	wire [31:0] r2243_out;
	wire [31:0] r2244_out;
	wire [31:0] r2245_out;
	wire [31:0] r2246_out;
	wire [31:0] r2247_out;
	wire [31:0] r2248_out;
	wire [31:0] r2249_out;
	wire [31:0] r2250_out;
	wire [31:0] r2251_out;
	wire [31:0] r2252_out;
	wire [31:0] r2253_out;
	wire [31:0] r2254_out;
	wire [31:0] r2255_out;
	wire [31:0] r2256_out;
	wire [31:0] r2257_out;
	wire [31:0] r2258_out;
	wire [31:0] r2259_out;
	wire [31:0] r2260_out;
	wire [31:0] r2261_out;
	wire [31:0] r2262_out;
	wire [31:0] r2263_out;
	wire [31:0] r2264_out;
	wire [31:0] r2265_out;
	wire [31:0] r2266_out;
	wire [31:0] r2267_out;
	wire [31:0] r2268_out;
	wire [31:0] r2269_out;
	wire [31:0] r2270_out;
	wire [31:0] r2271_out;
	wire [31:0] r2272_out;
	wire [31:0] r2273_out;
	wire [31:0] r2274_out;
	wire [31:0] r2275_out;
	wire [31:0] r2276_out;
	wire [31:0] r2277_out;
	wire [31:0] r2278_out;
	wire [31:0] r2279_out;
	wire [31:0] r2280_out;
	wire [31:0] r2281_out;
	wire [31:0] r2282_out;
	wire [31:0] r2283_out;
	wire [31:0] r2284_out;
	wire [31:0] r2285_out;
	wire [31:0] r2286_out;
	wire [31:0] r2287_out;
	wire [31:0] r2288_out;
	wire [31:0] r2289_out;
	wire [31:0] r2290_out;
	wire [31:0] r2291_out;
	wire [31:0] r2292_out;
	wire [31:0] r2293_out;
	wire [31:0] r2294_out;
	wire [31:0] r2295_out;
	wire [31:0] r2296_out;
	wire [31:0] r2297_out;
	wire [31:0] r2298_out;
	wire [31:0] r2299_out;
	wire [31:0] r2300_out;
	wire [31:0] r2301_out;
	wire [31:0] r2302_out;
	wire [31:0] r2303_out;
	wire [31:0] r2304_out;
	wire [31:0] r2305_out;
	wire [31:0] r2306_out;
	wire [31:0] r2307_out;
	wire [31:0] r2308_out;
	wire [31:0] r2309_out;
	wire [31:0] r2310_out;
	wire [31:0] r2311_out;
	wire [31:0] r2312_out;
	wire [31:0] r2313_out;
	wire [31:0] r2314_out;
	wire [31:0] r2315_out;
	wire [31:0] r2316_out;
	wire [31:0] r2317_out;
	wire [31:0] r2318_out;
	wire [31:0] r2319_out;
	wire [31:0] r2320_out;
	wire [31:0] r2321_out;
	wire [31:0] r2322_out;
	wire [31:0] r2323_out;
	wire [31:0] r2324_out;
	wire [31:0] r2325_out;
	wire [31:0] r2326_out;
	wire [31:0] r2327_out;
	wire [31:0] r2328_out;
	wire [31:0] r2329_out;
	wire [31:0] r2330_out;
	wire [31:0] r2331_out;
	wire [31:0] r2332_out;
	wire [31:0] r2333_out;
	wire [31:0] r2334_out;
	wire [31:0] r2335_out;
	wire [31:0] r2336_out;
	wire [31:0] r2337_out;
	wire [31:0] r2338_out;
	wire [31:0] r2339_out;
	wire [31:0] r2340_out;
	wire [31:0] r2341_out;
	wire [31:0] r2342_out;
	wire [31:0] r2343_out;
	wire [31:0] r2344_out;
	wire [31:0] r2345_out;
	wire [31:0] r2346_out;
	wire [31:0] r2347_out;
	wire [31:0] r2348_out;
	wire [31:0] r2349_out;
	wire [31:0] r2350_out;
	wire [31:0] r2351_out;
	wire [31:0] r2352_out;
	wire [31:0] r2353_out;
	wire [31:0] r2354_out;
	wire [31:0] r2355_out;
	wire [31:0] r2356_out;
	wire [31:0] r2357_out;
	wire [31:0] r2358_out;
	wire [31:0] r2359_out;
	wire [31:0] r2360_out;
	wire [31:0] r2361_out;
	wire [31:0] r2362_out;
	wire [31:0] r2363_out;
	wire [31:0] r2364_out;
	wire [31:0] r2365_out;
	wire [31:0] r2366_out;
	wire [31:0] r2367_out;
	wire [31:0] r2368_out;
	wire [31:0] r2369_out;
	wire [31:0] r2370_out;
	wire [31:0] r2371_out;
	wire [31:0] r2372_out;
	wire [31:0] r2373_out;
	wire [31:0] r2374_out;
	wire [31:0] r2375_out;
	wire [31:0] r2376_out;
	wire [31:0] r2377_out;
	wire [31:0] r2378_out;
	wire [31:0] r2379_out;
	wire [31:0] r2380_out;
	wire [31:0] r2381_out;
	wire [31:0] r2382_out;
	wire [31:0] r2383_out;
	wire [31:0] r2384_out;
	wire [31:0] r2385_out;
	wire [31:0] r2386_out;
	wire [31:0] r2387_out;
	wire [31:0] r2388_out;
	wire [31:0] r2389_out;
	wire [31:0] r2390_out;
	wire [31:0] r2391_out;
	wire [31:0] r2392_out;
	wire [31:0] r2393_out;
	wire [31:0] r2394_out;
	wire [31:0] r2395_out;
	wire [31:0] r2396_out;
	wire [31:0] r2397_out;
	wire [31:0] r2398_out;
	wire [31:0] r2399_out;
	wire [31:0] r2400_out;
	wire [31:0] r2401_out;
	wire [31:0] r2402_out;
	wire [31:0] r2403_out;
	wire [31:0] r2404_out;
	wire [31:0] r2405_out;
	wire [31:0] r2406_out;
	wire [31:0] r2407_out;
	wire [31:0] r2408_out;
	wire [31:0] r2409_out;
	wire [31:0] r2410_out;
	wire [31:0] r2411_out;
	wire [31:0] r2412_out;
	wire [31:0] r2413_out;
	wire [31:0] r2414_out;
	wire [31:0] r2415_out;
	wire [31:0] r2416_out;
	wire [31:0] r2417_out;
	wire [31:0] r2418_out;
	wire [31:0] r2419_out;
	wire [31:0] r2420_out;
	wire [31:0] r2421_out;
	wire [31:0] r2422_out;
	wire [31:0] r2423_out;
	wire [31:0] r2424_out;
	wire [31:0] r2425_out;
	wire [31:0] r2426_out;
	wire [31:0] r2427_out;
	wire [31:0] r2428_out;
	wire [31:0] r2429_out;
	wire [31:0] r2430_out;
	wire [31:0] r2431_out;
	wire [31:0] r2432_out;
	wire [31:0] r2433_out;
	wire [31:0] r2434_out;
	wire [31:0] r2435_out;
	wire [31:0] r2436_out;
	wire [31:0] r2437_out;
	wire [31:0] r2438_out;
	wire [31:0] r2439_out;
	wire [31:0] r2440_out;
	wire [31:0] r2441_out;
	wire [31:0] r2442_out;
	wire [31:0] r2443_out;
	wire [31:0] r2444_out;
	wire [31:0] r2445_out;
	wire [31:0] r2446_out;
	wire [31:0] r2447_out;
	wire [31:0] r2448_out;
	wire [31:0] r2449_out;
	wire [31:0] r2450_out;
	wire [31:0] r2451_out;
	wire [31:0] r2452_out;
	wire [31:0] r2453_out;
	wire [31:0] r2454_out;
	wire [31:0] r2455_out;
	wire [31:0] r2456_out;
	wire [31:0] r2457_out;
	wire [31:0] r2458_out;
	wire [31:0] r2459_out;
	wire [31:0] r2460_out;
	wire [31:0] r2461_out;
	wire [31:0] r2462_out;
	wire [31:0] r2463_out;
	wire [31:0] r2464_out;
	wire [31:0] r2465_out;
	wire [31:0] r2466_out;
	wire [31:0] r2467_out;
	wire [31:0] r2468_out;
	wire [31:0] r2469_out;
	wire [31:0] r2470_out;
	wire [31:0] r2471_out;
	wire [31:0] r2472_out;
	wire [31:0] r2473_out;
	wire [31:0] r2474_out;
	wire [31:0] r2475_out;
	wire [31:0] r2476_out;
	wire [31:0] r2477_out;
	wire [31:0] r2478_out;
	wire [31:0] r2479_out;
	wire [31:0] r2480_out;
	wire [31:0] r2481_out;
	wire [31:0] r2482_out;
	wire [31:0] r2483_out;
	wire [31:0] r2484_out;
	wire [31:0] r2485_out;
	wire [31:0] r2486_out;
	wire [31:0] r2487_out;
	wire [31:0] r2488_out;
	wire [31:0] r2489_out;
	wire [31:0] r2490_out;
	wire [31:0] r2491_out;
	wire [31:0] r2492_out;
	wire [31:0] r2493_out;
	wire [31:0] r2494_out;
	wire [31:0] r2495_out;
	wire [31:0] r2496_out;
	wire [31:0] r2497_out;
	wire [31:0] r2498_out;
	wire [31:0] r2499_out;
	wire [31:0] r2500_out;
	wire [31:0] r2501_out;
	wire [31:0] r2502_out;
	wire [31:0] r2503_out;
	wire [31:0] r2504_out;
	wire [31:0] r2505_out;
	wire [31:0] r2506_out;
	wire [31:0] r2507_out;
	wire [31:0] r2508_out;
	wire [31:0] r2509_out;
	wire [31:0] r2510_out;
	wire [31:0] r2511_out;
	wire [31:0] r2512_out;
	wire [31:0] r2513_out;
	wire [31:0] r2514_out;
	wire [31:0] r2515_out;
	wire [31:0] r2516_out;
	wire [31:0] r2517_out;
	wire [31:0] r2518_out;
	wire [31:0] r2519_out;
	wire [31:0] r2520_out;
	wire [31:0] r2521_out;
	wire [31:0] r2522_out;
	wire [31:0] r2523_out;
	wire [31:0] r2524_out;
	wire [31:0] r2525_out;
	wire [31:0] r2526_out;
	wire [31:0] r2527_out;
	wire [31:0] r2528_out;
	wire [31:0] r2529_out;
	wire [31:0] r2530_out;
	wire [31:0] r2531_out;
	wire [31:0] r2532_out;
	wire [31:0] r2533_out;
	wire [31:0] r2534_out;
	wire [31:0] r2535_out;
	wire [31:0] r2536_out;
	wire [31:0] r2537_out;
	wire [31:0] r2538_out;
	wire [31:0] r2539_out;
	wire [31:0] r2540_out;
	wire [31:0] r2541_out;
	wire [31:0] r2542_out;
	wire [31:0] r2543_out;
	wire [31:0] r2544_out;
	wire [31:0] r2545_out;
	wire [31:0] r2546_out;
	wire [31:0] r2547_out;
	wire [31:0] r2548_out;
	wire [31:0] r2549_out;
	wire [31:0] r2550_out;
	wire [31:0] r2551_out;
	wire [31:0] r2552_out;
	wire [31:0] r2553_out;
	wire [31:0] r2554_out;
	wire [31:0] r2555_out;
	wire [31:0] r2556_out;
	wire [31:0] r2557_out;
	wire [31:0] r2558_out;
	wire [31:0] r2559_out;
	wire [31:0] r2560_out;
	wire [31:0] r2561_out;
	wire [31:0] r2562_out;
	wire [31:0] r2563_out;
	wire [31:0] r2564_out;
	wire [31:0] r2565_out;
	wire [31:0] r2566_out;
	wire [31:0] r2567_out;
	wire [31:0] r2568_out;
	wire [31:0] r2569_out;
	wire [31:0] r2570_out;
	wire [31:0] r2571_out;
	wire [31:0] r2572_out;
	wire [31:0] r2573_out;
	wire [31:0] r2574_out;
	wire [31:0] r2575_out;
	wire [31:0] r2576_out;
	wire [31:0] r2577_out;
	wire [31:0] r2578_out;
	wire [31:0] r2579_out;
	wire [31:0] r2580_out;
	wire [31:0] r2581_out;
	wire [31:0] r2582_out;
	wire [31:0] r2583_out;
	wire [31:0] r2584_out;
	wire [31:0] r2585_out;
	wire [31:0] r2586_out;
	wire [31:0] r2587_out;
	wire [31:0] r2588_out;
	wire [31:0] r2589_out;
	wire [31:0] r2590_out;
	wire [31:0] r2591_out;
	wire [31:0] r2592_out;
	wire [31:0] r2593_out;
	wire [31:0] r2594_out;
	wire [31:0] r2595_out;
	wire [31:0] r2596_out;
	wire [31:0] r2597_out;
	wire [31:0] r2598_out;
	wire [31:0] r2599_out;
	wire [31:0] r2600_out;
	wire [31:0] r2601_out;
	wire [31:0] r2602_out;
	wire [31:0] r2603_out;
	wire [31:0] r2604_out;
	wire [31:0] r2605_out;
	wire [31:0] r2606_out;
	wire [31:0] r2607_out;
	wire [31:0] r2608_out;
	wire [31:0] r2609_out;
	wire [31:0] r2610_out;
	wire [31:0] r2611_out;
	wire [31:0] r2612_out;
	wire [31:0] r2613_out;
	wire [31:0] r2614_out;
	wire [31:0] r2615_out;
	wire [31:0] r2616_out;
	wire [31:0] r2617_out;
	wire [31:0] r2618_out;
	wire [31:0] r2619_out;
	wire [31:0] r2620_out;
	wire [31:0] r2621_out;
	wire [31:0] r2622_out;
	wire [31:0] r2623_out;
	wire [31:0] r2624_out;
	wire [31:0] r2625_out;
	wire [31:0] r2626_out;
	wire [31:0] r2627_out;
	wire [31:0] r2628_out;
	wire [31:0] r2629_out;
	wire [31:0] r2630_out;
	wire [31:0] r2631_out;
	wire [31:0] r2632_out;
	wire [31:0] r2633_out;
	wire [31:0] r2634_out;
	wire [31:0] r2635_out;
	wire [31:0] r2636_out;
	wire [31:0] r2637_out;
	wire [31:0] r2638_out;
	wire [31:0] r2639_out;
	wire [31:0] r2640_out;
	wire [31:0] r2641_out;
	wire [31:0] r2642_out;
	wire [31:0] r2643_out;
	wire [31:0] r2644_out;
	wire [31:0] r2645_out;
	wire [31:0] r2646_out;
	wire [31:0] r2647_out;
	wire [31:0] r2648_out;
	wire [31:0] r2649_out;
	wire [31:0] r2650_out;
	wire [31:0] r2651_out;
	wire [31:0] r2652_out;
	wire [31:0] r2653_out;
	wire [31:0] r2654_out;
	wire [31:0] r2655_out;
	wire [31:0] r2656_out;
	wire [31:0] r2657_out;
	wire [31:0] r2658_out;
	wire [31:0] r2659_out;
	wire [31:0] r2660_out;
	wire [31:0] r2661_out;
	wire [31:0] r2662_out;
	wire [31:0] r2663_out;
	wire [31:0] r2664_out;
	wire [31:0] r2665_out;
	wire [31:0] r2666_out;
	wire [31:0] r2667_out;
	wire [31:0] r2668_out;
	wire [31:0] r2669_out;
	wire [31:0] r2670_out;
	wire [31:0] r2671_out;
	wire [31:0] r2672_out;
	wire [31:0] r2673_out;
	wire [31:0] r2674_out;
	wire [31:0] r2675_out;
	wire [31:0] r2676_out;
	wire [31:0] r2677_out;
	wire [31:0] r2678_out;
	wire [31:0] r2679_out;
	wire [31:0] r2680_out;
	wire [31:0] r2681_out;
	wire [31:0] r2682_out;
	wire [31:0] r2683_out;
	wire [31:0] r2684_out;
	wire [31:0] r2685_out;
	wire [31:0] r2686_out;
	wire [31:0] r2687_out;
	wire [31:0] r2688_out;
	wire [31:0] r2689_out;
	wire [31:0] r2690_out;
	wire [31:0] r2691_out;
	wire [31:0] r2692_out;
	wire [31:0] r2693_out;
	wire [31:0] r2694_out;
	wire [31:0] r2695_out;
	wire [31:0] r2696_out;
	wire [31:0] r2697_out;
	wire [31:0] r2698_out;
	wire [31:0] r2699_out;
	wire [31:0] r2700_out;
	wire [31:0] r2701_out;
	wire [31:0] r2702_out;
	wire [31:0] r2703_out;
	wire [31:0] r2704_out;
	wire [31:0] r2705_out;
	wire [31:0] r2706_out;
	wire [31:0] r2707_out;
	wire [31:0] r2708_out;
	wire [31:0] r2709_out;
	wire [31:0] r2710_out;
	wire [31:0] r2711_out;
	wire [31:0] r2712_out;
	wire [31:0] r2713_out;
	wire [31:0] r2714_out;
	wire [31:0] r2715_out;
	wire [31:0] r2716_out;
	wire [31:0] r2717_out;
	wire [31:0] r2718_out;
	wire [31:0] r2719_out;
	wire [31:0] r2720_out;
	wire [31:0] r2721_out;
	wire [31:0] r2722_out;
	wire [31:0] r2723_out;
	wire [31:0] r2724_out;
	wire [31:0] r2725_out;
	wire [31:0] r2726_out;
	wire [31:0] r2727_out;
	wire [31:0] r2728_out;
	wire [31:0] r2729_out;
	wire [31:0] r2730_out;
	wire [31:0] r2731_out;
	wire [31:0] r2732_out;
	wire [31:0] r2733_out;
	wire [31:0] r2734_out;
	wire [31:0] r2735_out;
	wire [31:0] r2736_out;
	wire [31:0] r2737_out;
	wire [31:0] r2738_out;
	wire [31:0] r2739_out;
	wire [31:0] r2740_out;
	wire [31:0] r2741_out;
	wire [31:0] r2742_out;
	wire [31:0] r2743_out;
	wire [31:0] r2744_out;
	wire [31:0] r2745_out;
	wire [31:0] r2746_out;
	wire [31:0] r2747_out;
	wire [31:0] r2748_out;
	wire [31:0] r2749_out;
	wire [31:0] r2750_out;
	wire [31:0] r2751_out;
	wire [31:0] r2752_out;
	wire [31:0] r2753_out;
	wire [31:0] r2754_out;
	wire [31:0] r2755_out;
	wire [31:0] r2756_out;
	wire [31:0] r2757_out;
	wire [31:0] r2758_out;
	wire [31:0] r2759_out;
	wire [31:0] r2760_out;
	wire [31:0] r2761_out;
	wire [31:0] r2762_out;
	wire [31:0] r2763_out;
	wire [31:0] r2764_out;
	wire [31:0] r2765_out;
	wire [31:0] r2766_out;
	wire [31:0] r2767_out;
	wire [31:0] r2768_out;
	wire [31:0] r2769_out;
	wire [31:0] r2770_out;
	wire [31:0] r2771_out;
	wire [31:0] r2772_out;
	wire [31:0] r2773_out;
	wire [31:0] r2774_out;
	wire [31:0] r2775_out;
	wire [31:0] r2776_out;
	wire [31:0] r2777_out;
	wire [31:0] r2778_out;
	wire [31:0] r2779_out;
	wire [31:0] r2780_out;
	wire [31:0] r2781_out;
	wire [31:0] r2782_out;
	wire [31:0] r2783_out;
	wire [31:0] r2784_out;
	wire [31:0] r2785_out;
	wire [31:0] r2786_out;
	wire [31:0] r2787_out;
	wire [31:0] r2788_out;
	wire [31:0] r2789_out;
	wire [31:0] r2790_out;
	wire [31:0] r2791_out;
	wire [31:0] r2792_out;
	wire [31:0] r2793_out;
	wire [31:0] r2794_out;
	wire [31:0] r2795_out;
	wire [31:0] r2796_out;
	wire [31:0] r2797_out;
	wire [31:0] r2798_out;
	wire [31:0] r2799_out;
	wire [31:0] r2800_out;
	wire [31:0] r2801_out;
	wire [31:0] r2802_out;
	wire [31:0] r2803_out;
	wire [31:0] r2804_out;
	wire [31:0] r2805_out;
	wire [31:0] r2806_out;
	wire [31:0] r2807_out;
	wire [31:0] r2808_out;
	wire [31:0] r2809_out;
	wire [31:0] r2810_out;
	wire [31:0] r2811_out;
	wire [31:0] r2812_out;
	wire [31:0] r2813_out;
	wire [31:0] r2814_out;
	wire [31:0] r2815_out;
	wire [31:0] r2816_out;
	wire [31:0] r2817_out;
	wire [31:0] r2818_out;
	wire [31:0] r2819_out;
	wire [31:0] r2820_out;
	wire [31:0] r2821_out;
	wire [31:0] r2822_out;
	wire [31:0] r2823_out;
	wire [31:0] r2824_out;
	wire [31:0] r2825_out;
	wire [31:0] r2826_out;
	wire [31:0] r2827_out;
	wire [31:0] r2828_out;
	wire [31:0] r2829_out;
	wire [31:0] r2830_out;
	wire [31:0] r2831_out;
	wire [31:0] r2832_out;
	wire [31:0] r2833_out;
	wire [31:0] r2834_out;
	wire [31:0] r2835_out;
	wire [31:0] r2836_out;
	wire [31:0] r2837_out;
	wire [31:0] r2838_out;
	wire [31:0] r2839_out;
	wire [31:0] r2840_out;
	wire [31:0] r2841_out;
	wire [31:0] r2842_out;
	wire [31:0] r2843_out;
	wire [31:0] r2844_out;
	wire [31:0] r2845_out;
	wire [31:0] r2846_out;
	wire [31:0] r2847_out;
	wire [31:0] r2848_out;
	wire [31:0] r2849_out;
	wire [31:0] r2850_out;
	wire [31:0] r2851_out;
	wire [31:0] r2852_out;
	wire [31:0] r2853_out;
	wire [31:0] r2854_out;
	wire [31:0] r2855_out;
	wire [31:0] r2856_out;
	wire [31:0] r2857_out;
	wire [31:0] r2858_out;
	wire [31:0] r2859_out;
	wire [31:0] r2860_out;
	wire [31:0] r2861_out;
	wire [31:0] r2862_out;
	wire [31:0] r2863_out;
	wire [31:0] r2864_out;
	wire [31:0] r2865_out;
	wire [31:0] r2866_out;
	wire [31:0] r2867_out;
	wire [31:0] r2868_out;
	wire [31:0] r2869_out;
	wire [31:0] r2870_out;
	wire [31:0] r2871_out;
	wire [31:0] r2872_out;
	wire [31:0] r2873_out;
	wire [31:0] r2874_out;
	wire [31:0] r2875_out;
	wire [31:0] r2876_out;
	wire [31:0] r2877_out;
	wire [31:0] r2878_out;
	wire [31:0] r2879_out;
	wire [31:0] r2880_out;
	wire [31:0] r2881_out;
	wire [31:0] r2882_out;
	wire [31:0] r2883_out;
	wire [31:0] r2884_out;
	wire [31:0] r2885_out;
	wire [31:0] r2886_out;
	wire [31:0] r2887_out;
	wire [31:0] r2888_out;
	wire [31:0] r2889_out;
	wire [31:0] r2890_out;
	wire [31:0] r2891_out;
	wire [31:0] r2892_out;
	wire [31:0] r2893_out;
	wire [31:0] r2894_out;
	wire [31:0] r2895_out;
	wire [31:0] r2896_out;
	wire [31:0] r2897_out;
	wire [31:0] r2898_out;
	wire [31:0] r2899_out;
	wire [31:0] r2900_out;
	wire [31:0] r2901_out;
	wire [31:0] r2902_out;
	wire [31:0] r2903_out;
	wire [31:0] r2904_out;
	wire [31:0] r2905_out;
	wire [31:0] r2906_out;
	wire [31:0] r2907_out;
	wire [31:0] r2908_out;
	wire [31:0] r2909_out;
	wire [31:0] r2910_out;
	wire [31:0] r2911_out;
	wire [31:0] r2912_out;
	wire [31:0] r2913_out;
	wire [31:0] r2914_out;
	wire [31:0] r2915_out;
	wire [31:0] r2916_out;
	wire [31:0] r2917_out;
	wire [31:0] r2918_out;
	wire [31:0] r2919_out;
	wire [31:0] r2920_out;
	wire [31:0] r2921_out;
	wire [31:0] r2922_out;
	wire [31:0] r2923_out;
	wire [31:0] r2924_out;
	wire [31:0] r2925_out;
	wire [31:0] r2926_out;
	wire [31:0] r2927_out;
	wire [31:0] r2928_out;
	wire [31:0] r2929_out;
	wire [31:0] r2930_out;
	wire [31:0] r2931_out;
	wire [31:0] r2932_out;
	wire [31:0] r2933_out;
	wire [31:0] r2934_out;
	wire [31:0] r2935_out;
	wire [31:0] r2936_out;
	wire [31:0] r2937_out;
	wire [31:0] r2938_out;
	wire [31:0] r2939_out;
	wire [31:0] r2940_out;
	wire [31:0] r2941_out;
	wire [31:0] r2942_out;
	wire [31:0] r2943_out;
	wire [31:0] r2944_out;
	wire [31:0] r2945_out;
	wire [31:0] r2946_out;
	wire [31:0] r2947_out;
	wire [31:0] r2948_out;
	wire [31:0] r2949_out;
	wire [31:0] r2950_out;
	wire [31:0] r2951_out;
	wire [31:0] r2952_out;
	wire [31:0] r2953_out;
	wire [31:0] r2954_out;
	wire [31:0] r2955_out;
	wire [31:0] r2956_out;
	wire [31:0] r2957_out;
	wire [31:0] r2958_out;
	wire [31:0] r2959_out;
	wire [31:0] r2960_out;
	wire [31:0] r2961_out;
	wire [31:0] r2962_out;
	wire [31:0] r2963_out;
	wire [31:0] r2964_out;
	wire [31:0] r2965_out;
	wire [31:0] r2966_out;
	wire [31:0] r2967_out;
	wire [31:0] r2968_out;
	wire [31:0] r2969_out;
	wire [31:0] r2970_out;
	wire [31:0] r2971_out;
	wire [31:0] r2972_out;
	wire [31:0] r2973_out;
	wire [31:0] r2974_out;
	wire [31:0] r2975_out;
	wire [31:0] r2976_out;
	wire [31:0] r2977_out;
	wire [31:0] r2978_out;
	wire [31:0] r2979_out;
	wire [31:0] r2980_out;
	wire [31:0] r2981_out;
	wire [31:0] r2982_out;
	wire [31:0] r2983_out;
	wire [31:0] r2984_out;
	wire [31:0] r2985_out;
	wire [31:0] r2986_out;
	wire [31:0] r2987_out;
	wire [31:0] r2988_out;
	wire [31:0] r2989_out;
	wire [31:0] r2990_out;
	wire [31:0] r2991_out;
	wire [31:0] r2992_out;
	wire [31:0] r2993_out;
	wire [31:0] r2994_out;
	wire [31:0] r2995_out;
	wire [31:0] r2996_out;
	wire [31:0] r2997_out;
	wire [31:0] r2998_out;
	wire [31:0] r2999_out;
	wire [31:0] r3000_out;
	wire [31:0] r3001_out;
	wire [31:0] r3002_out;
	wire [31:0] r3003_out;
	wire [31:0] r3004_out;
	wire [31:0] r3005_out;
	wire [31:0] r3006_out;
	wire [31:0] r3007_out;
	wire [31:0] r3008_out;
	wire [31:0] r3009_out;
	wire [31:0] r3010_out;
	wire [31:0] r3011_out;
	wire [31:0] r3012_out;
	wire [31:0] r3013_out;
	wire [31:0] r3014_out;
	wire [31:0] r3015_out;
	wire [31:0] r3016_out;
	wire [31:0] r3017_out;
	wire [31:0] r3018_out;
	wire [31:0] r3019_out;
	wire [31:0] r3020_out;
	wire [31:0] r3021_out;
	wire [31:0] r3022_out;
	wire [31:0] r3023_out;
	wire [31:0] r3024_out;
	wire [31:0] r3025_out;
	wire [31:0] r3026_out;
	wire [31:0] r3027_out;
	wire [31:0] r3028_out;
	wire [31:0] r3029_out;
	wire [31:0] r3030_out;
	wire [31:0] r3031_out;
	wire [31:0] r3032_out;
	wire [31:0] r3033_out;
	wire [31:0] r3034_out;
	wire [31:0] r3035_out;
	wire [31:0] r3036_out;
	wire [31:0] r3037_out;
	wire [31:0] r3038_out;
	wire [31:0] r3039_out;
	wire [31:0] r3040_out;
	wire [31:0] r3041_out;
	wire [31:0] r3042_out;
	wire [31:0] r3043_out;
	wire [31:0] r3044_out;
	wire [31:0] r3045_out;
	wire [31:0] r3046_out;
	wire [31:0] r3047_out;
	wire [31:0] r3048_out;
	wire [31:0] r3049_out;
	wire [31:0] r3050_out;
	wire [31:0] r3051_out;
	wire [31:0] r3052_out;
	wire [31:0] r3053_out;
	wire [31:0] r3054_out;
	wire [31:0] r3055_out;
	wire [31:0] r3056_out;
	wire [31:0] r3057_out;
	wire [31:0] r3058_out;
	wire [31:0] r3059_out;
	wire [31:0] r3060_out;
	wire [31:0] r3061_out;
	wire [31:0] r3062_out;
	wire [31:0] r3063_out;
	wire [31:0] r3064_out;
	wire [31:0] r3065_out;
	wire [31:0] r3066_out;
	wire [31:0] r3067_out;
	wire [31:0] r3068_out;
	wire [31:0] r3069_out;
	wire [31:0] r3070_out;
	wire [31:0] r3071_out;
	wire [31:0] r3072_out;
	wire [31:0] r3073_out;
	wire [31:0] r3074_out;
	wire [31:0] r3075_out;
	wire [31:0] r3076_out;
	wire [31:0] r3077_out;
	wire [31:0] r3078_out;
	wire [31:0] r3079_out;
	wire [31:0] r3080_out;
	wire [31:0] r3081_out;
	wire [31:0] r3082_out;
	wire [31:0] r3083_out;
	wire [31:0] r3084_out;
	wire [31:0] r3085_out;
	wire [31:0] r3086_out;
	wire [31:0] r3087_out;
	wire [31:0] r3088_out;
	wire [31:0] r3089_out;
	wire [31:0] r3090_out;
	wire [31:0] r3091_out;
	wire [31:0] r3092_out;
	wire [31:0] r3093_out;
	wire [31:0] r3094_out;
	wire [31:0] r3095_out;
	wire [31:0] r3096_out;
	wire [31:0] r3097_out;
	wire [31:0] r3098_out;
	wire [31:0] r3099_out;
	wire [31:0] r3100_out;
	wire [31:0] r3101_out;
	wire [31:0] r3102_out;
	wire [31:0] r3103_out;
	wire [31:0] r3104_out;
	wire [31:0] r3105_out;
	wire [31:0] r3106_out;
	wire [31:0] r3107_out;
	wire [31:0] r3108_out;
	wire [31:0] r3109_out;
	wire [31:0] r3110_out;
	wire [31:0] r3111_out;
	wire [31:0] r3112_out;
	wire [31:0] r3113_out;
	wire [31:0] r3114_out;
	wire [31:0] r3115_out;
	wire [31:0] r3116_out;
	wire [31:0] r3117_out;
	wire [31:0] r3118_out;
	wire [31:0] r3119_out;
	wire [31:0] r3120_out;
	wire [31:0] r3121_out;
	wire [31:0] r3122_out;
	wire [31:0] r3123_out;
	wire [31:0] r3124_out;
	wire [31:0] r3125_out;
	wire [31:0] r3126_out;
	wire [31:0] r3127_out;
	wire [31:0] r3128_out;
	wire [31:0] r3129_out;
	wire [31:0] r3130_out;
	wire [31:0] r3131_out;
	wire [31:0] r3132_out;
	wire [31:0] r3133_out;
	wire [31:0] r3134_out;
	wire [31:0] r3135_out;
	wire [31:0] r3136_out;
	wire [31:0] r3137_out;
	wire [31:0] r3138_out;
	wire [31:0] r3139_out;
	wire [31:0] r3140_out;
	wire [31:0] r3141_out;
	wire [31:0] r3142_out;
	wire [31:0] r3143_out;
	wire [31:0] r3144_out;
	wire [31:0] r3145_out;
	wire [31:0] r3146_out;
	wire [31:0] r3147_out;
	wire [31:0] r3148_out;
	wire [31:0] r3149_out;
	wire [31:0] r3150_out;
	wire [31:0] r3151_out;
	wire [31:0] r3152_out;
	wire [31:0] r3153_out;
	wire [31:0] r3154_out;
	wire [31:0] r3155_out;
	wire [31:0] r3156_out;
	wire [31:0] r3157_out;
	wire [31:0] r3158_out;
	wire [31:0] r3159_out;
	wire [31:0] r3160_out;
	wire [31:0] r3161_out;
	wire [31:0] r3162_out;
	wire [31:0] r3163_out;
	wire [31:0] r3164_out;
	wire [31:0] r3165_out;
	wire [31:0] r3166_out;
	wire [31:0] r3167_out;
	wire [31:0] r3168_out;
	wire [31:0] r3169_out;
	wire [31:0] r3170_out;
	wire [31:0] r3171_out;
	wire [31:0] r3172_out;
	wire [31:0] r3173_out;
	wire [31:0] r3174_out;
	wire [31:0] r3175_out;
	wire [31:0] r3176_out;
	wire [31:0] r3177_out;
	wire [31:0] r3178_out;
	wire [31:0] r3179_out;
	wire [31:0] r3180_out;
	wire [31:0] r3181_out;
	wire [31:0] r3182_out;
	wire [31:0] r3183_out;
	wire [31:0] r3184_out;
	wire [31:0] r3185_out;
	wire [31:0] r3186_out;
	wire [31:0] r3187_out;
	wire [31:0] r3188_out;
	wire [31:0] r3189_out;
	wire [31:0] r3190_out;
	wire [31:0] r3191_out;
	wire [31:0] r3192_out;
	wire [31:0] r3193_out;
	wire [31:0] r3194_out;
	wire [31:0] r3195_out;
	wire [31:0] r3196_out;
	wire [31:0] r3197_out;
	wire [31:0] r3198_out;
	wire [31:0] r3199_out;
	wire [31:0] r3200_out;
	wire [31:0] r3201_out;
	wire [31:0] r3202_out;
	wire [31:0] r3203_out;
	wire [31:0] r3204_out;
	wire [31:0] r3205_out;
	wire [31:0] r3206_out;
	wire [31:0] r3207_out;
	wire [31:0] r3208_out;
	wire [31:0] r3209_out;
	wire [31:0] r3210_out;
	wire [31:0] r3211_out;
	wire [31:0] r3212_out;
	wire [31:0] r3213_out;
	wire [31:0] r3214_out;
	wire [31:0] r3215_out;
	wire [31:0] r3216_out;
	wire [31:0] r3217_out;
	wire [31:0] r3218_out;
	wire [31:0] r3219_out;
	wire [31:0] r3220_out;
	wire [31:0] r3221_out;
	wire [31:0] r3222_out;
	wire [31:0] r3223_out;
	wire [31:0] r3224_out;
	wire [31:0] r3225_out;
	wire [31:0] r3226_out;
	wire [31:0] r3227_out;
	wire [31:0] r3228_out;
	wire [31:0] r3229_out;
	wire [31:0] r3230_out;
	wire [31:0] r3231_out;
	wire [31:0] r3232_out;
	wire [31:0] r3233_out;
	wire [31:0] r3234_out;
	wire [31:0] r3235_out;
	wire [31:0] r3236_out;
	wire [31:0] r3237_out;
	wire [31:0] r3238_out;
	wire [31:0] r3239_out;
	wire [31:0] r3240_out;
	wire [31:0] r3241_out;
	wire [31:0] r3242_out;
	wire [31:0] r3243_out;
	wire [31:0] r3244_out;
	wire [31:0] r3245_out;
	wire [31:0] r3246_out;
	wire [31:0] r3247_out;
	wire [31:0] r3248_out;
	wire [31:0] r3249_out;
	wire [31:0] r3250_out;
	wire [31:0] r3251_out;
	wire [31:0] r3252_out;
	wire [31:0] r3253_out;
	wire [31:0] r3254_out;
	wire [31:0] r3255_out;
	wire [31:0] r3256_out;
	wire [31:0] r3257_out;
	wire [31:0] r3258_out;
	wire [31:0] r3259_out;
	wire [31:0] r3260_out;
	wire [31:0] r3261_out;
	wire [31:0] r3262_out;
	wire [31:0] r3263_out;
	wire [31:0] r3264_out;
	wire [31:0] r3265_out;
	wire [31:0] r3266_out;
	wire [31:0] r3267_out;
	wire [31:0] r3268_out;
	wire [31:0] r3269_out;
	wire [31:0] r3270_out;
	wire [31:0] r3271_out;
	wire [31:0] r3272_out;
	wire [31:0] r3273_out;
	wire [31:0] r3274_out;
	wire [31:0] r3275_out;
	wire [31:0] r3276_out;
	wire [31:0] r3277_out;
	wire [31:0] r3278_out;
	wire [31:0] r3279_out;
	wire [31:0] r3280_out;
	wire [31:0] r3281_out;
	wire [31:0] r3282_out;
	wire [31:0] r3283_out;
	wire [31:0] r3284_out;
	wire [31:0] r3285_out;
	wire [31:0] r3286_out;
	wire [31:0] r3287_out;
	wire [31:0] r3288_out;
	wire [31:0] r3289_out;
	wire [31:0] r3290_out;
	wire [31:0] r3291_out;
	wire [31:0] r3292_out;
	wire [31:0] r3293_out;
	wire [31:0] r3294_out;
	wire [31:0] r3295_out;
	wire [31:0] r3296_out;
	wire [31:0] r3297_out;
	wire [31:0] r3298_out;
	wire [31:0] r3299_out;
	wire [31:0] r3300_out;
	wire [31:0] r3301_out;
	wire [31:0] r3302_out;
	wire [31:0] r3303_out;
	wire [31:0] r3304_out;
	wire [31:0] r3305_out;
	wire [31:0] r3306_out;
	wire [31:0] r3307_out;
	wire [31:0] r3308_out;
	wire [31:0] r3309_out;
	wire [31:0] r3310_out;
	wire [31:0] r3311_out;
	wire [31:0] r3312_out;
	wire [31:0] r3313_out;
	wire [31:0] r3314_out;
	wire [31:0] r3315_out;
	wire [31:0] r3316_out;
	wire [31:0] r3317_out;
	wire [31:0] r3318_out;
	wire [31:0] r3319_out;
	wire [31:0] r3320_out;
	wire [31:0] r3321_out;
	wire [31:0] r3322_out;
	wire [31:0] r3323_out;
	wire [31:0] r3324_out;
	wire [31:0] r3325_out;
	wire [31:0] r3326_out;
	wire [31:0] r3327_out;
	wire [31:0] r3328_out;
	wire [31:0] r3329_out;
	wire [31:0] r3330_out;
	wire [31:0] r3331_out;
	wire [31:0] r3332_out;
	wire [31:0] r3333_out;
	wire [31:0] r3334_out;
	wire [31:0] r3335_out;
	wire [31:0] r3336_out;
	wire [31:0] r3337_out;
	wire [31:0] r3338_out;
	wire [31:0] r3339_out;
	wire [31:0] r3340_out;
	wire [31:0] r3341_out;
	wire [31:0] r3342_out;
	wire [31:0] r3343_out;
	wire [31:0] r3344_out;
	wire [31:0] r3345_out;
	wire [31:0] r3346_out;
	wire [31:0] r3347_out;
	wire [31:0] r3348_out;
	wire [31:0] r3349_out;
	wire [31:0] r3350_out;
	wire [31:0] r3351_out;
	wire [31:0] r3352_out;
	wire [31:0] r3353_out;
	wire [31:0] r3354_out;
	wire [31:0] r3355_out;
	wire [31:0] r3356_out;
	wire [31:0] r3357_out;
	wire [31:0] r3358_out;
	wire [31:0] r3359_out;
	wire [31:0] r3360_out;
	wire [31:0] r3361_out;
	wire [31:0] r3362_out;
	wire [31:0] r3363_out;
	wire [31:0] r3364_out;
	wire [31:0] r3365_out;
	wire [31:0] r3366_out;
	wire [31:0] r3367_out;
	wire [31:0] r3368_out;
	wire [31:0] r3369_out;
	wire [31:0] r3370_out;
	wire [31:0] r3371_out;
	wire [31:0] r3372_out;
	wire [31:0] r3373_out;
	wire [31:0] r3374_out;
	wire [31:0] r3375_out;
	wire [31:0] r3376_out;
	wire [31:0] r3377_out;
	wire [31:0] r3378_out;
	wire [31:0] r3379_out;
	wire [31:0] r3380_out;
	wire [31:0] r3381_out;
	wire [31:0] r3382_out;
	wire [31:0] r3383_out;
	wire [31:0] r3384_out;
	wire [31:0] r3385_out;
	wire [31:0] r3386_out;
	wire [31:0] r3387_out;
	wire [31:0] r3388_out;
	wire [31:0] r3389_out;
	wire [31:0] r3390_out;
	wire [31:0] r3391_out;
	wire [31:0] r3392_out;
	wire [31:0] r3393_out;
	wire [31:0] r3394_out;
	wire [31:0] r3395_out;
	wire [31:0] r3396_out;
	wire [31:0] r3397_out;
	wire [31:0] r3398_out;
	wire [31:0] r3399_out;
	wire [31:0] r3400_out;
	wire [31:0] r3401_out;
	wire [31:0] r3402_out;
	wire [31:0] r3403_out;
	wire [31:0] r3404_out;
	wire [31:0] r3405_out;
	wire [31:0] r3406_out;
	wire [31:0] r3407_out;
	wire [31:0] r3408_out;
	wire [31:0] r3409_out;
	wire [31:0] r3410_out;
	wire [31:0] r3411_out;
	wire [31:0] r3412_out;
	wire [31:0] r3413_out;
	wire [31:0] r3414_out;
	wire [31:0] r3415_out;
	wire [31:0] r3416_out;
	wire [31:0] r3417_out;
	wire [31:0] r3418_out;
	wire [31:0] r3419_out;
	wire [31:0] r3420_out;
	wire [31:0] r3421_out;
	wire [31:0] r3422_out;
	wire [31:0] r3423_out;
	wire [31:0] r3424_out;
	wire [31:0] r3425_out;
	wire [31:0] r3426_out;
	wire [31:0] r3427_out;
	wire [31:0] r3428_out;
	wire [31:0] r3429_out;
	wire [31:0] r3430_out;
	wire [31:0] r3431_out;
	wire [31:0] r3432_out;
	wire [31:0] r3433_out;
	wire [31:0] r3434_out;
	wire [31:0] r3435_out;
	wire [31:0] r3436_out;
	wire [31:0] r3437_out;
	wire [31:0] r3438_out;
	wire [31:0] r3439_out;
	wire [31:0] r3440_out;
	wire [31:0] r3441_out;
	wire [31:0] r3442_out;
	wire [31:0] r3443_out;
	wire [31:0] r3444_out;
	wire [31:0] r3445_out;
	wire [31:0] r3446_out;
	wire [31:0] r3447_out;
	wire [31:0] r3448_out;
	wire [31:0] r3449_out;
	wire [31:0] r3450_out;
	wire [31:0] r3451_out;
	wire [31:0] r3452_out;
	wire [31:0] r3453_out;
	wire [31:0] r3454_out;
	wire [31:0] r3455_out;
	wire [31:0] r3456_out;
	wire [31:0] r3457_out;
	wire [31:0] r3458_out;
	wire [31:0] r3459_out;
	wire [31:0] r3460_out;
	wire [31:0] r3461_out;
	wire [31:0] r3462_out;
	wire [31:0] r3463_out;
	wire [31:0] r3464_out;
	wire [31:0] r3465_out;
	wire [31:0] r3466_out;
	wire [31:0] r3467_out;
	wire [31:0] r3468_out;
	wire [31:0] r3469_out;
	wire [31:0] r3470_out;
	wire [31:0] r3471_out;
	wire [31:0] r3472_out;
	wire [31:0] r3473_out;
	wire [31:0] r3474_out;
	wire [31:0] r3475_out;
	wire [31:0] r3476_out;
	wire [31:0] r3477_out;
	wire [31:0] r3478_out;
	wire [31:0] r3479_out;
	wire [31:0] r3480_out;
	wire [31:0] r3481_out;
	wire [31:0] r3482_out;
	wire [31:0] r3483_out;
	wire [31:0] r3484_out;
	wire [31:0] r3485_out;
	wire [31:0] r3486_out;
	wire [31:0] r3487_out;
	wire [31:0] r3488_out;
	wire [31:0] r3489_out;
	wire [31:0] r3490_out;
	wire [31:0] r3491_out;
	wire [31:0] r3492_out;
	wire [31:0] r3493_out;
	wire [31:0] r3494_out;
	wire [31:0] r3495_out;
	wire [31:0] r3496_out;
	wire [31:0] r3497_out;
	wire [31:0] r3498_out;
	wire [31:0] r3499_out;
	wire [31:0] r3500_out;
	wire [31:0] r3501_out;
	wire [31:0] r3502_out;
	wire [31:0] r3503_out;
	wire [31:0] r3504_out;
	wire [31:0] r3505_out;
	wire [31:0] r3506_out;
	wire [31:0] r3507_out;
	wire [31:0] r3508_out;
	wire [31:0] r3509_out;
	wire [31:0] r3510_out;
	wire [31:0] r3511_out;
	wire [31:0] r3512_out;
	wire [31:0] r3513_out;
	wire [31:0] r3514_out;
	wire [31:0] r3515_out;
	wire [31:0] r3516_out;
	wire [31:0] r3517_out;
	wire [31:0] r3518_out;
	wire [31:0] r3519_out;
	wire [31:0] r3520_out;
	wire [31:0] r3521_out;
	wire [31:0] r3522_out;
	wire [31:0] r3523_out;
	wire [31:0] r3524_out;
	wire [31:0] r3525_out;
	wire [31:0] r3526_out;
	wire [31:0] r3527_out;
	wire [31:0] r3528_out;
	wire [31:0] r3529_out;
	wire [31:0] r3530_out;
	wire [31:0] r3531_out;
	wire [31:0] r3532_out;
	wire [31:0] r3533_out;
	wire [31:0] r3534_out;
	wire [31:0] r3535_out;
	wire [31:0] r3536_out;
	wire [31:0] r3537_out;
	wire [31:0] r3538_out;
	wire [31:0] r3539_out;
	wire [31:0] r3540_out;
	wire [31:0] r3541_out;
	wire [31:0] r3542_out;
	wire [31:0] r3543_out;
	wire [31:0] r3544_out;
	wire [31:0] r3545_out;
	wire [31:0] r3546_out;
	wire [31:0] r3547_out;
	wire [31:0] r3548_out;
	wire [31:0] r3549_out;
	wire [31:0] r3550_out;
	wire [31:0] r3551_out;
	wire [31:0] r3552_out;
	wire [31:0] r3553_out;
	wire [31:0] r3554_out;
	wire [31:0] r3555_out;
	wire [31:0] r3556_out;
	wire [31:0] r3557_out;
	wire [31:0] r3558_out;
	wire [31:0] r3559_out;
	wire [31:0] r3560_out;
	wire [31:0] r3561_out;
	wire [31:0] r3562_out;
	wire [31:0] r3563_out;
	wire [31:0] r3564_out;
	wire [31:0] r3565_out;
	wire [31:0] r3566_out;
	wire [31:0] r3567_out;
	wire [31:0] r3568_out;
	wire [31:0] r3569_out;
	wire [31:0] r3570_out;
	wire [31:0] r3571_out;
	wire [31:0] r3572_out;
	wire [31:0] r3573_out;
	wire [31:0] r3574_out;
	wire [31:0] r3575_out;
	wire [31:0] r3576_out;
	wire [31:0] r3577_out;
	wire [31:0] r3578_out;
	wire [31:0] r3579_out;
	wire [31:0] r3580_out;
	wire [31:0] r3581_out;
	wire [31:0] r3582_out;
	wire [31:0] r3583_out;
	wire [31:0] r3584_out;
	wire [31:0] r3585_out;
	wire [31:0] r3586_out;
	wire [31:0] r3587_out;
	wire [31:0] r3588_out;
	wire [31:0] r3589_out;
	wire [31:0] r3590_out;
	wire [31:0] r3591_out;
	wire [31:0] r3592_out;
	wire [31:0] r3593_out;
	wire [31:0] r3594_out;
	wire [31:0] r3595_out;
	wire [31:0] r3596_out;
	wire [31:0] r3597_out;
	wire [31:0] r3598_out;
	wire [31:0] r3599_out;
	wire [31:0] r3600_out;
	wire [31:0] r3601_out;
	wire [31:0] r3602_out;
	wire [31:0] r3603_out;
	wire [31:0] r3604_out;
	wire [31:0] r3605_out;
	wire [31:0] r3606_out;
	wire [31:0] r3607_out;
	wire [31:0] r3608_out;
	wire [31:0] r3609_out;
	wire [31:0] r3610_out;
	wire [31:0] r3611_out;
	wire [31:0] r3612_out;
	wire [31:0] r3613_out;
	wire [31:0] r3614_out;
	wire [31:0] r3615_out;
	wire [31:0] r3616_out;
	wire [31:0] r3617_out;
	wire [31:0] r3618_out;
	wire [31:0] r3619_out;
	wire [31:0] r3620_out;
	wire [31:0] r3621_out;
	wire [31:0] r3622_out;
	wire [31:0] r3623_out;
	wire [31:0] r3624_out;
	wire [31:0] r3625_out;
	wire [31:0] r3626_out;
	wire [31:0] r3627_out;
	wire [31:0] r3628_out;
	wire [31:0] r3629_out;
	wire [31:0] r3630_out;
	wire [31:0] r3631_out;
	wire [31:0] r3632_out;
	wire [31:0] r3633_out;
	wire [31:0] r3634_out;
	wire [31:0] r3635_out;
	wire [31:0] r3636_out;
	wire [31:0] r3637_out;
	wire [31:0] r3638_out;
	wire [31:0] r3639_out;
	wire [31:0] r3640_out;
	wire [31:0] r3641_out;
	wire [31:0] r3642_out;
	wire [31:0] r3643_out;
	wire [31:0] r3644_out;
	wire [31:0] r3645_out;
	wire [31:0] r3646_out;
	wire [31:0] r3647_out;
	wire [31:0] r3648_out;
	wire [31:0] r3649_out;
	wire [31:0] r3650_out;
	wire [31:0] r3651_out;
	wire [31:0] r3652_out;
	wire [31:0] r3653_out;
	wire [31:0] r3654_out;
	wire [31:0] r3655_out;
	wire [31:0] r3656_out;
	wire [31:0] r3657_out;
	wire [31:0] r3658_out;
	wire [31:0] r3659_out;
	wire [31:0] r3660_out;
	wire [31:0] r3661_out;
	wire [31:0] r3662_out;
	wire [31:0] r3663_out;
	wire [31:0] r3664_out;
	wire [31:0] r3665_out;
	wire [31:0] r3666_out;
	wire [31:0] r3667_out;
	wire [31:0] r3668_out;
	wire [31:0] r3669_out;
	wire [31:0] r3670_out;
	wire [31:0] r3671_out;
	wire [31:0] r3672_out;
	wire [31:0] r3673_out;
	wire [31:0] r3674_out;
	wire [31:0] r3675_out;
	wire [31:0] r3676_out;
	wire [31:0] r3677_out;
	wire [31:0] r3678_out;
	wire [31:0] r3679_out;
	wire [31:0] r3680_out;
	wire [31:0] r3681_out;
	wire [31:0] r3682_out;
	wire [31:0] r3683_out;
	wire [31:0] r3684_out;
	wire [31:0] r3685_out;
	wire [31:0] r3686_out;
	wire [31:0] r3687_out;
	wire [31:0] r3688_out;
	wire [31:0] r3689_out;
	wire [31:0] r3690_out;
	wire [31:0] r3691_out;
	wire [31:0] r3692_out;
	wire [31:0] r3693_out;
	wire [31:0] r3694_out;
	wire [31:0] r3695_out;
	wire [31:0] r3696_out;
	wire [31:0] r3697_out;
	wire [31:0] r3698_out;
	wire [31:0] r3699_out;
	wire [31:0] r3700_out;
	wire [31:0] r3701_out;
	wire [31:0] r3702_out;
	wire [31:0] r3703_out;
	wire [31:0] r3704_out;
	wire [31:0] r3705_out;
	wire [31:0] r3706_out;
	wire [31:0] r3707_out;
	wire [31:0] r3708_out;
	wire [31:0] r3709_out;
	wire [31:0] r3710_out;
	wire [31:0] r3711_out;
	wire [31:0] r3712_out;
	wire [31:0] r3713_out;
	wire [31:0] r3714_out;
	wire [31:0] r3715_out;
	wire [31:0] r3716_out;
	wire [31:0] r3717_out;
	wire [31:0] r3718_out;
	wire [31:0] r3719_out;
	wire [31:0] r3720_out;
	wire [31:0] r3721_out;
	wire [31:0] r3722_out;
	wire [31:0] r3723_out;
	wire [31:0] r3724_out;
	wire [31:0] r3725_out;
	wire [31:0] r3726_out;
	wire [31:0] r3727_out;
	wire [31:0] r3728_out;
	wire [31:0] r3729_out;
	wire [31:0] r3730_out;
	wire [31:0] r3731_out;
	wire [31:0] r3732_out;
	wire [31:0] r3733_out;
	wire [31:0] r3734_out;
	wire [31:0] r3735_out;
	wire [31:0] r3736_out;
	wire [31:0] r3737_out;
	wire [31:0] r3738_out;
	wire [31:0] r3739_out;
	wire [31:0] r3740_out;
	wire [31:0] r3741_out;
	wire [31:0] r3742_out;
	wire [31:0] r3743_out;
	wire [31:0] r3744_out;
	wire [31:0] r3745_out;
	wire [31:0] r3746_out;
	wire [31:0] r3747_out;
	wire [31:0] r3748_out;
	wire [31:0] r3749_out;
	wire [31:0] r3750_out;
	wire [31:0] r3751_out;
	wire [31:0] r3752_out;
	wire [31:0] r3753_out;
	wire [31:0] r3754_out;
	wire [31:0] r3755_out;
	wire [31:0] r3756_out;
	wire [31:0] r3757_out;
	wire [31:0] r3758_out;
	wire [31:0] r3759_out;
	wire [31:0] r3760_out;
	wire [31:0] r3761_out;
	wire [31:0] r3762_out;
	wire [31:0] r3763_out;
	wire [31:0] r3764_out;
	wire [31:0] r3765_out;
	wire [31:0] r3766_out;
	wire [31:0] r3767_out;
	wire [31:0] r3768_out;
	wire [31:0] r3769_out;
	wire [31:0] r3770_out;
	wire [31:0] r3771_out;
	wire [31:0] r3772_out;
	wire [31:0] r3773_out;
	wire [31:0] r3774_out;
	wire [31:0] r3775_out;
	wire [31:0] r3776_out;
	wire [31:0] r3777_out;
	wire [31:0] r3778_out;
	wire [31:0] r3779_out;
	wire [31:0] r3780_out;
	wire [31:0] r3781_out;
	wire [31:0] r3782_out;
	wire [31:0] r3783_out;
	wire [31:0] r3784_out;
	wire [31:0] r3785_out;
	wire [31:0] r3786_out;
	wire [31:0] r3787_out;
	wire [31:0] r3788_out;
	wire [31:0] r3789_out;
	wire [31:0] r3790_out;
	wire [31:0] r3791_out;
	wire [31:0] r3792_out;
	wire [31:0] r3793_out;
	wire [31:0] r3794_out;
	wire [31:0] r3795_out;
	wire [31:0] r3796_out;
	wire [31:0] r3797_out;
	wire [31:0] r3798_out;
	wire [31:0] r3799_out;
	wire [31:0] r3800_out;
	wire [31:0] r3801_out;
	wire [31:0] r3802_out;
	wire [31:0] r3803_out;
	wire [31:0] r3804_out;
	wire [31:0] r3805_out;
	wire [31:0] r3806_out;
	wire [31:0] r3807_out;
	wire [31:0] r3808_out;
	wire [31:0] r3809_out;
	wire [31:0] r3810_out;
	wire [31:0] r3811_out;
	wire [31:0] r3812_out;
	wire [31:0] r3813_out;
	wire [31:0] r3814_out;
	wire [31:0] r3815_out;
	wire [31:0] r3816_out;
	wire [31:0] r3817_out;
	wire [31:0] r3818_out;
	wire [31:0] r3819_out;
	wire [31:0] r3820_out;
	wire [31:0] r3821_out;
	wire [31:0] r3822_out;
	wire [31:0] r3823_out;
	wire [31:0] r3824_out;
	wire [31:0] r3825_out;
	wire [31:0] r3826_out;
	wire [31:0] r3827_out;
	wire [31:0] r3828_out;
	wire [31:0] r3829_out;
	wire [31:0] r3830_out;
	wire [31:0] r3831_out;
	wire [31:0] r3832_out;
	wire [31:0] r3833_out;
	wire [31:0] r3834_out;
	wire [31:0] r3835_out;
	wire [31:0] r3836_out;
	wire [31:0] r3837_out;
	wire [31:0] r3838_out;
	wire [31:0] r3839_out;
	wire [31:0] r3840_out;
	wire [31:0] r3841_out;
	wire [31:0] r3842_out;
	wire [31:0] r3843_out;
	wire [31:0] r3844_out;
	wire [31:0] r3845_out;
	wire [31:0] r3846_out;
	wire [31:0] r3847_out;
	wire [31:0] r3848_out;
	wire [31:0] r3849_out;
	wire [31:0] r3850_out;
	wire [31:0] r3851_out;
	wire [31:0] r3852_out;
	wire [31:0] r3853_out;
	wire [31:0] r3854_out;
	wire [31:0] r3855_out;
	wire [31:0] r3856_out;
	wire [31:0] r3857_out;
	wire [31:0] r3858_out;
	wire [31:0] r3859_out;
	wire [31:0] r3860_out;
	wire [31:0] r3861_out;
	wire [31:0] r3862_out;
	wire [31:0] r3863_out;
	wire [31:0] r3864_out;
	wire [31:0] r3865_out;
	wire [31:0] r3866_out;
	wire [31:0] r3867_out;
	wire [31:0] r3868_out;
	wire [31:0] r3869_out;
	wire [31:0] r3870_out;
	wire [31:0] r3871_out;
	wire [31:0] r3872_out;
	wire [31:0] r3873_out;
	wire [31:0] r3874_out;
	wire [31:0] r3875_out;
	wire [31:0] r3876_out;
	wire [31:0] r3877_out;
	wire [31:0] r3878_out;
	wire [31:0] r3879_out;
	wire [31:0] r3880_out;
	wire [31:0] r3881_out;
	wire [31:0] r3882_out;
	wire [31:0] r3883_out;
	wire [31:0] r3884_out;
	wire [31:0] r3885_out;
	wire [31:0] r3886_out;
	wire [31:0] r3887_out;
	wire [31:0] r3888_out;
	wire [31:0] r3889_out;
	wire [31:0] r3890_out;
	wire [31:0] r3891_out;
	wire [31:0] r3892_out;
	wire [31:0] r3893_out;
	wire [31:0] r3894_out;
	wire [31:0] r3895_out;
	wire [31:0] r3896_out;
	wire [31:0] r3897_out;
	wire [31:0] r3898_out;
	wire [31:0] r3899_out;
	wire [31:0] r3900_out;
	wire [31:0] r3901_out;
	wire [31:0] r3902_out;
	wire [31:0] r3903_out;
	wire [31:0] r3904_out;
	wire [31:0] r3905_out;
	wire [31:0] r3906_out;
	wire [31:0] r3907_out;
	wire [31:0] r3908_out;
	wire [31:0] r3909_out;
	wire [31:0] r3910_out;
	wire [31:0] r3911_out;
	wire [31:0] r3912_out;
	wire [31:0] r3913_out;
	wire [31:0] r3914_out;
	wire [31:0] r3915_out;
	wire [31:0] r3916_out;
	wire [31:0] r3917_out;
	wire [31:0] r3918_out;
	wire [31:0] r3919_out;
	wire [31:0] r3920_out;
	wire [31:0] r3921_out;
	wire [31:0] r3922_out;
	wire [31:0] r3923_out;
	wire [31:0] r3924_out;
	wire [31:0] r3925_out;
	wire [31:0] r3926_out;
	wire [31:0] r3927_out;
	wire [31:0] r3928_out;
	wire [31:0] r3929_out;
	wire [31:0] r3930_out;
	wire [31:0] r3931_out;
	wire [31:0] r3932_out;
	wire [31:0] r3933_out;
	wire [31:0] r3934_out;
	wire [31:0] r3935_out;
	wire [31:0] r3936_out;
	wire [31:0] r3937_out;
	wire [31:0] r3938_out;
	wire [31:0] r3939_out;
	wire [31:0] r3940_out;
	wire [31:0] r3941_out;
	wire [31:0] r3942_out;
	wire [31:0] r3943_out;
	wire [31:0] r3944_out;
	wire [31:0] r3945_out;
	wire [31:0] r3946_out;
	wire [31:0] r3947_out;
	wire [31:0] r3948_out;
	wire [31:0] r3949_out;
	wire [31:0] r3950_out;
	wire [31:0] r3951_out;
	wire [31:0] r3952_out;
	wire [31:0] r3953_out;
	wire [31:0] r3954_out;
	wire [31:0] r3955_out;
	wire [31:0] r3956_out;
	wire [31:0] r3957_out;
	wire [31:0] r3958_out;
	wire [31:0] r3959_out;
	wire [31:0] r3960_out;
	wire [31:0] r3961_out;
	wire [31:0] r3962_out;
	wire [31:0] r3963_out;
	wire [31:0] r3964_out;
	wire [31:0] r3965_out;
	wire [31:0] r3966_out;
	wire [31:0] r3967_out;
	wire [31:0] r3968_out;
	wire [31:0] r3969_out;
	wire [31:0] r3970_out;
	wire [31:0] r3971_out;
	wire [31:0] r3972_out;
	wire [31:0] r3973_out;
	wire [31:0] r3974_out;
	wire [31:0] r3975_out;
	wire [31:0] r3976_out;
	wire [31:0] r3977_out;
	wire [31:0] r3978_out;
	wire [31:0] r3979_out;
	wire [31:0] r3980_out;
	wire [31:0] r3981_out;
	wire [31:0] r3982_out;
	wire [31:0] r3983_out;
	wire [31:0] r3984_out;
	wire [31:0] r3985_out;
	wire [31:0] r3986_out;
	wire [31:0] r3987_out;
	wire [31:0] r3988_out;
	wire [31:0] r3989_out;
	wire [31:0] r3990_out;
	wire [31:0] r3991_out;
	wire [31:0] r3992_out;
	wire [31:0] r3993_out;
	wire [31:0] r3994_out;
	wire [31:0] r3995_out;
	wire [31:0] r3996_out;
	wire [31:0] r3997_out;
	wire [31:0] r3998_out;
	wire [31:0] r3999_out;
	wire [31:0] r4000_out;
	wire [31:0] r4001_out;
	wire [31:0] r4002_out;
	wire [31:0] r4003_out;
	wire [31:0] r4004_out;
	wire [31:0] r4005_out;
	wire [31:0] r4006_out;
	wire [31:0] r4007_out;
	wire [31:0] r4008_out;
	wire [31:0] r4009_out;
	wire [31:0] r4010_out;
	wire [31:0] r4011_out;
	wire [31:0] r4012_out;
	wire [31:0] r4013_out;
	wire [31:0] r4014_out;
	wire [31:0] r4015_out;
	wire [31:0] r4016_out;
	wire [31:0] r4017_out;
	wire [31:0] r4018_out;
	wire [31:0] r4019_out;
	wire [31:0] r4020_out;
	wire [31:0] r4021_out;
	wire [31:0] r4022_out;
	wire [31:0] r4023_out;
	wire [31:0] r4024_out;
	wire [31:0] r4025_out;
	wire [31:0] r4026_out;
	wire [31:0] r4027_out;
	wire [31:0] r4028_out;
	wire [31:0] r4029_out;
	wire [31:0] r4030_out;
	wire [31:0] r4031_out;
	wire [31:0] r4032_out;
	wire [31:0] r4033_out;
	wire [31:0] r4034_out;
	wire [31:0] r4035_out;
	wire [31:0] r4036_out;
	wire [31:0] r4037_out;
	wire [31:0] r4038_out;
	wire [31:0] r4039_out;
	wire [31:0] r4040_out;
	wire [31:0] r4041_out;
	wire [31:0] r4042_out;
	wire [31:0] r4043_out;
	wire [31:0] r4044_out;
	wire [31:0] r4045_out;
	wire [31:0] r4046_out;
	wire [31:0] r4047_out;
	wire [31:0] r4048_out;
	wire [31:0] r4049_out;
	wire [31:0] r4050_out;
	wire [31:0] r4051_out;
	wire [31:0] r4052_out;
	wire [31:0] r4053_out;
	wire [31:0] r4054_out;
	wire [31:0] r4055_out;
	wire [31:0] r4056_out;
	wire [31:0] r4057_out;
	wire [31:0] r4058_out;
	wire [31:0] r4059_out;
	wire [31:0] r4060_out;
	wire [31:0] r4061_out;
	wire [31:0] r4062_out;
	wire [31:0] r4063_out;
	wire [31:0] r4064_out;
	wire [31:0] r4065_out;
	wire [31:0] r4066_out;
	wire [31:0] r4067_out;
	wire [31:0] r4068_out;
	wire [31:0] r4069_out;
	wire [31:0] r4070_out;
	wire [31:0] r4071_out;
	wire [31:0] r4072_out;
	wire [31:0] r4073_out;
	wire [31:0] r4074_out;
	wire [31:0] r4075_out;
	wire [31:0] r4076_out;
	wire [31:0] r4077_out;
	wire [31:0] r4078_out;
	wire [31:0] r4079_out;
	wire [31:0] r4080_out;
	wire [31:0] r4081_out;
	wire [31:0] r4082_out;
	wire [31:0] r4083_out;
	wire [31:0] r4084_out;
	wire [31:0] r4085_out;
	wire [31:0] r4086_out;
	wire [31:0] r4087_out;
	wire [31:0] r4088_out;
	wire [31:0] r4089_out;
	wire [31:0] r4090_out;
	wire [31:0] r4091_out;
	wire [31:0] r4092_out;
	wire [31:0] r4093_out;
	wire [31:0] r4094_out;
	wire [31:0] r4095_out;
	wire [31:0] r4096_out;
	wire [31:0] r4097_out;
	wire [31:0] r4098_out;
	wire [31:0] r4099_out;
	wire [31:0] r4100_out;
	wire [31:0] r4101_out;
	wire [31:0] r4102_out;
	wire [31:0] r4103_out;
	wire [31:0] r4104_out;
	wire [31:0] r4105_out;
	wire [31:0] r4106_out;
	wire [31:0] r4107_out;
	wire [31:0] r4108_out;
	wire [31:0] r4109_out;
	wire [31:0] r4110_out;
	wire [31:0] r4111_out;
	wire [31:0] r4112_out;
	wire [31:0] r4113_out;
	wire [31:0] r4114_out;
	wire [31:0] r4115_out;
	wire [31:0] r4116_out;
	wire [31:0] r4117_out;
	wire [31:0] r4118_out;
	wire [31:0] r4119_out;
	wire [31:0] r4120_out;
	wire [31:0] r4121_out;
	wire [31:0] r4122_out;
	wire [31:0] r4123_out;
	wire [31:0] r4124_out;
	wire [31:0] r4125_out;
	wire [31:0] r4126_out;
	wire [31:0] r4127_out;
	wire [31:0] r4128_out;
	wire [31:0] r4129_out;
	wire [31:0] r4130_out;
	wire [31:0] r4131_out;
	wire [31:0] r4132_out;
	wire [31:0] r4133_out;
	wire [31:0] r4134_out;
	wire [31:0] r4135_out;
	wire [31:0] r4136_out;
	wire [31:0] r4137_out;
	wire [31:0] r4138_out;
	wire [31:0] r4139_out;
	wire [31:0] r4140_out;
	wire [31:0] r4141_out;
	wire [31:0] r4142_out;
	wire [31:0] r4143_out;
	wire [31:0] r4144_out;
	wire [31:0] r4145_out;
	wire [31:0] r4146_out;
	wire [31:0] r4147_out;
	wire [31:0] r4148_out;
	wire [31:0] r4149_out;
	wire [31:0] r4150_out;
	wire [31:0] r4151_out;
	wire [31:0] r4152_out;
	wire [31:0] r4153_out;
	wire [31:0] r4154_out;
	wire [31:0] r4155_out;
	wire [31:0] r4156_out;
	wire [31:0] r4157_out;
	wire [31:0] r4158_out;
	wire [31:0] r4159_out;
	wire [31:0] r4160_out;
	wire [31:0] r4161_out;
	wire [31:0] r4162_out;
	wire [31:0] r4163_out;
	wire [31:0] r4164_out;
	wire [31:0] r4165_out;
	wire [31:0] r4166_out;
	wire [31:0] r4167_out;
	wire [31:0] r4168_out;
	wire [31:0] r4169_out;
	wire [31:0] r4170_out;
	wire [31:0] r4171_out;
	wire [31:0] r4172_out;
	wire [31:0] r4173_out;
	wire [31:0] r4174_out;
	wire [31:0] r4175_out;
	wire [31:0] r4176_out;
	wire [31:0] r4177_out;
	wire [31:0] r4178_out;
	wire [31:0] r4179_out;
	wire [31:0] r4180_out;
	wire [31:0] r4181_out;
	wire [31:0] r4182_out;
	wire [31:0] r4183_out;
	wire [31:0] r4184_out;
	wire [31:0] r4185_out;
	wire [31:0] r4186_out;
	wire [31:0] r4187_out;
	wire [31:0] r4188_out;
	wire [31:0] r4189_out;
	wire [31:0] r4190_out;
	wire [31:0] r4191_out;
	wire [31:0] r4192_out;
	wire [31:0] r4193_out;
	wire [31:0] r4194_out;
	wire [31:0] r4195_out;
	wire [31:0] r4196_out;
	wire [31:0] r4197_out;
	wire [31:0] r4198_out;
	wire [31:0] r4199_out;
	wire [31:0] r4200_out;
	wire [31:0] r4201_out;
	wire [31:0] r4202_out;
	wire [31:0] r4203_out;
	wire [31:0] r4204_out;
	wire [31:0] r4205_out;
	wire [31:0] r4206_out;
	wire [31:0] r4207_out;
	wire [31:0] r4208_out;
	wire [31:0] r4209_out;
	wire [31:0] r4210_out;
	wire [31:0] r4211_out;
	wire [31:0] r4212_out;
	wire [31:0] r4213_out;
	wire [31:0] r4214_out;
	wire [31:0] r4215_out;
	wire [31:0] r4216_out;
	wire [31:0] r4217_out;
	wire [31:0] r4218_out;
	wire [31:0] r4219_out;
	wire [31:0] r4220_out;
	wire [31:0] r4221_out;
	wire [31:0] r4222_out;
	wire [31:0] r4223_out;
	wire [31:0] r4224_out;
	wire [31:0] r4225_out;
	wire [31:0] r4226_out;
	wire [31:0] r4227_out;
	wire [31:0] r4228_out;
	wire [31:0] r4229_out;
	wire [31:0] r4230_out;
	wire [31:0] r4231_out;
	wire [31:0] r4232_out;
	wire [31:0] r4233_out;
	wire [31:0] r4234_out;
	wire [31:0] r4235_out;
	wire [31:0] r4236_out;
	wire [31:0] r4237_out;
	wire [31:0] r4238_out;
	wire [31:0] r4239_out;
	wire [31:0] r4240_out;
	wire [31:0] r4241_out;
	wire [31:0] r4242_out;
	wire [31:0] r4243_out;
	wire [31:0] r4244_out;
	wire [31:0] r4245_out;
	wire [31:0] r4246_out;
	wire [31:0] r4247_out;
	wire [31:0] r4248_out;
	wire [31:0] r4249_out;
	wire [31:0] r4250_out;
	wire [31:0] r4251_out;
	wire [31:0] r4252_out;
	wire [31:0] r4253_out;
	wire [31:0] r4254_out;
	wire [31:0] r4255_out;
	wire [31:0] r4256_out;
	wire [31:0] r4257_out;
	wire [31:0] r4258_out;
	wire [31:0] r4259_out;
	wire [31:0] r4260_out;
	wire [31:0] r4261_out;
	wire [31:0] r4262_out;
	wire [31:0] r4263_out;
	wire [31:0] r4264_out;
	wire [31:0] r4265_out;
	wire [31:0] r4266_out;
	wire [31:0] r4267_out;
	wire [31:0] r4268_out;
	wire [31:0] r4269_out;
	wire [31:0] r4270_out;
	wire [31:0] r4271_out;
	wire [31:0] r4272_out;
	wire [31:0] r4273_out;
	wire [31:0] r4274_out;
	wire [31:0] r4275_out;
	wire [31:0] r4276_out;
	wire [31:0] r4277_out;
	wire [31:0] r4278_out;
	wire [31:0] r4279_out;
	wire [31:0] r4280_out;
	wire [31:0] r4281_out;
	wire [31:0] r4282_out;
	wire [31:0] r4283_out;
	wire [31:0] r4284_out;
	wire [31:0] r4285_out;
	wire [31:0] r4286_out;
	wire [31:0] r4287_out;
	wire [31:0] r4288_out;
	wire [31:0] r4289_out;
	wire [31:0] r4290_out;
	wire [31:0] r4291_out;
	wire [31:0] r4292_out;
	wire [31:0] r4293_out;
	wire [31:0] r4294_out;
	wire [31:0] r4295_out;
	wire [31:0] r4296_out;
	wire [31:0] r4297_out;
	wire [31:0] r4298_out;
	wire [31:0] r4299_out;
	wire [31:0] r4300_out;
	wire [31:0] r4301_out;
	wire [31:0] r4302_out;
	wire [31:0] r4303_out;
	wire [31:0] r4304_out;
	wire [31:0] r4305_out;
	wire [31:0] r4306_out;
	wire [31:0] r4307_out;
	wire [31:0] r4308_out;
	wire [31:0] r4309_out;
	wire [31:0] r4310_out;
	wire [31:0] r4311_out;
	wire [31:0] r4312_out;
	wire [31:0] r4313_out;
	wire [31:0] r4314_out;
	wire [31:0] r4315_out;
	wire [31:0] r4316_out;
	wire [31:0] r4317_out;
	wire [31:0] r4318_out;
	wire [31:0] r4319_out;
	wire [31:0] r4320_out;
	wire [31:0] r4321_out;
	wire [31:0] r4322_out;
	wire [31:0] r4323_out;
	wire [31:0] r4324_out;
	wire [31:0] r4325_out;
	wire [31:0] r4326_out;
	wire [31:0] r4327_out;
	wire [31:0] r4328_out;
	wire [31:0] r4329_out;
	wire [31:0] r4330_out;
	wire [31:0] r4331_out;
	wire [31:0] r4332_out;
	wire [31:0] r4333_out;
	wire [31:0] r4334_out;
	wire [31:0] r4335_out;
	wire [31:0] r4336_out;
	wire [31:0] r4337_out;
	wire [31:0] r4338_out;
	wire [31:0] r4339_out;
	wire [31:0] r4340_out;
	wire [31:0] r4341_out;
	wire [31:0] r4342_out;
	wire [31:0] r4343_out;
	wire [31:0] r4344_out;
	wire [31:0] r4345_out;
	wire [31:0] r4346_out;
	wire [31:0] r4347_out;
	wire [31:0] r4348_out;
	wire [31:0] r4349_out;
	wire [31:0] r4350_out;
	wire [31:0] r4351_out;
	wire [31:0] r4352_out;
	wire [31:0] r4353_out;
	wire [31:0] r4354_out;
	wire [31:0] r4355_out;
	wire [31:0] r4356_out;
	wire [31:0] r4357_out;
	wire [31:0] r4358_out;
	wire [31:0] r4359_out;
	wire [31:0] r4360_out;
	wire [31:0] r4361_out;
	wire [31:0] r4362_out;
	wire [31:0] r4363_out;
	wire [31:0] r4364_out;
	wire [31:0] r4365_out;
	wire [31:0] r4366_out;
	wire [31:0] r4367_out;
	wire [31:0] r4368_out;
	wire [31:0] r4369_out;
	wire [31:0] r4370_out;
	wire [31:0] r4371_out;
	wire [31:0] r4372_out;
	wire [31:0] r4373_out;
	wire [31:0] r4374_out;
	wire [31:0] r4375_out;
	wire [31:0] r4376_out;
	wire [31:0] r4377_out;
	wire [31:0] r4378_out;
	wire [31:0] r4379_out;
	wire [31:0] r4380_out;
	wire [31:0] r4381_out;
	wire [31:0] r4382_out;
	wire [31:0] r4383_out;
	wire [31:0] r4384_out;
	wire [31:0] r4385_out;
	wire [31:0] r4386_out;
	wire [31:0] r4387_out;
	wire [31:0] r4388_out;
	wire [31:0] r4389_out;
	wire [31:0] r4390_out;
	wire [31:0] r4391_out;
	wire [31:0] r4392_out;
	wire [31:0] r4393_out;
	wire [31:0] r4394_out;
	wire [31:0] r4395_out;
	wire [31:0] r4396_out;
	wire [31:0] r4397_out;
	wire [31:0] r4398_out;
	wire [31:0] r4399_out;
	wire [31:0] r4400_out;
	wire [31:0] r4401_out;
	wire [31:0] r4402_out;
	wire [31:0] r4403_out;
	wire [31:0] r4404_out;
	wire [31:0] r4405_out;
	wire [31:0] r4406_out;
	wire [31:0] r4407_out;
	wire [31:0] r4408_out;
	wire [31:0] r4409_out;
	wire [31:0] r4410_out;
	wire [31:0] r4411_out;
	wire [31:0] r4412_out;
	wire [31:0] r4413_out;
	wire [31:0] r4414_out;
	wire [31:0] r4415_out;
	wire [31:0] r4416_out;
	wire [31:0] r4417_out;
	wire [31:0] r4418_out;
	wire [31:0] r4419_out;
	wire [31:0] r4420_out;
	wire [31:0] r4421_out;
	wire [31:0] r4422_out;
	wire [31:0] r4423_out;
	wire [31:0] r4424_out;
	wire [31:0] r4425_out;
	wire [31:0] r4426_out;
	wire [31:0] r4427_out;
	wire [31:0] r4428_out;
	wire [31:0] r4429_out;
	wire [31:0] r4430_out;
	wire [31:0] r4431_out;
	wire [31:0] r4432_out;
	wire [31:0] r4433_out;
	wire [31:0] r4434_out;
	wire [31:0] r4435_out;
	wire [31:0] r4436_out;
	wire [31:0] r4437_out;
	wire [31:0] r4438_out;
	wire [31:0] r4439_out;
	wire [31:0] r4440_out;
	wire [31:0] r4441_out;
	wire [31:0] r4442_out;
	wire [31:0] r4443_out;
	wire [31:0] r4444_out;
	wire [31:0] r4445_out;
	wire [31:0] r4446_out;
	wire [31:0] r4447_out;
	wire [31:0] r4448_out;
	wire [31:0] r4449_out;
	wire [31:0] r4450_out;
	wire [31:0] r4451_out;
	wire [31:0] r4452_out;
	wire [31:0] r4453_out;
	wire [31:0] r4454_out;
	wire [31:0] r4455_out;
	wire [31:0] r4456_out;
	wire [31:0] r4457_out;
	wire [31:0] r4458_out;
	wire [31:0] r4459_out;
	wire [31:0] r4460_out;
	wire [31:0] r4461_out;
	wire [31:0] r4462_out;
	wire [31:0] r4463_out;
	wire [31:0] r4464_out;
	wire [31:0] r4465_out;
	wire [31:0] r4466_out;
	wire [31:0] r4467_out;
	wire [31:0] r4468_out;
	wire [31:0] r4469_out;
	wire [31:0] r4470_out;
	wire [31:0] r4471_out;
	wire [31:0] r4472_out;
	wire [31:0] r4473_out;
	wire [31:0] r4474_out;
	wire [31:0] r4475_out;
	wire [31:0] r4476_out;
	wire [31:0] r4477_out;
	wire [31:0] r4478_out;
	wire [31:0] r4479_out;
	wire [31:0] r4480_out;
	wire [31:0] r4481_out;
	wire [31:0] r4482_out;
	wire [31:0] r4483_out;
	wire [31:0] r4484_out;
	wire [31:0] r4485_out;
	wire [31:0] r4486_out;
	wire [31:0] r4487_out;
	wire [31:0] r4488_out;
	wire [31:0] r4489_out;
	wire [31:0] r4490_out;
	wire [31:0] r4491_out;
	wire [31:0] r4492_out;
	wire [31:0] r4493_out;
	wire [31:0] r4494_out;
	wire [31:0] r4495_out;
	wire [31:0] r4496_out;
	wire [31:0] r4497_out;
	wire [31:0] r4498_out;
	wire [31:0] r4499_out;
	wire [31:0] r4500_out;
	wire [31:0] r4501_out;
	wire [31:0] r4502_out;
	wire [31:0] r4503_out;
	wire [31:0] r4504_out;
	wire [31:0] r4505_out;
	wire [31:0] r4506_out;
	wire [31:0] r4507_out;
	wire [31:0] r4508_out;
	wire [31:0] r4509_out;
	wire [31:0] r4510_out;
	wire [31:0] r4511_out;
	wire [31:0] r4512_out;
	wire [31:0] r4513_out;
	wire [31:0] r4514_out;
	wire [31:0] r4515_out;
	wire [31:0] r4516_out;
	wire [31:0] r4517_out;
	wire [31:0] r4518_out;
	wire [31:0] r4519_out;
	wire [31:0] r4520_out;
	wire [31:0] r4521_out;
	wire [31:0] r4522_out;
	wire [31:0] r4523_out;
	wire [31:0] r4524_out;
	wire [31:0] r4525_out;
	wire [31:0] r4526_out;
	wire [31:0] r4527_out;
	wire [31:0] r4528_out;
	wire [31:0] r4529_out;
	wire [31:0] r4530_out;
	wire [31:0] r4531_out;
	wire [31:0] r4532_out;
	wire [31:0] r4533_out;
	wire [31:0] r4534_out;
	wire [31:0] r4535_out;
	wire [31:0] r4536_out;
	wire [31:0] r4537_out;
	wire [31:0] r4538_out;
	wire [31:0] r4539_out;
	wire [31:0] r4540_out;
	wire [31:0] r4541_out;
	wire [31:0] r4542_out;
	wire [31:0] r4543_out;
	wire [31:0] r4544_out;
	wire [31:0] r4545_out;
	wire [31:0] r4546_out;
	wire [31:0] r4547_out;
	wire [31:0] r4548_out;
	wire [31:0] r4549_out;
	wire [31:0] r4550_out;
	wire [31:0] r4551_out;
	wire [31:0] r4552_out;
	wire [31:0] r4553_out;
	wire [31:0] r4554_out;
	wire [31:0] r4555_out;
	wire [31:0] r4556_out;
	wire [31:0] r4557_out;
	wire [31:0] r4558_out;
	wire [31:0] r4559_out;
	wire [31:0] r4560_out;
	wire [31:0] r4561_out;
	wire [31:0] r4562_out;
	wire [31:0] r4563_out;
	wire [31:0] r4564_out;
	wire [31:0] r4565_out;
	wire [31:0] r4566_out;
	wire [31:0] r4567_out;
	wire [31:0] r4568_out;
	wire [31:0] r4569_out;
	wire [31:0] r4570_out;
	wire [31:0] r4571_out;
	wire [31:0] r4572_out;
	wire [31:0] r4573_out;
	wire [31:0] r4574_out;
	wire [31:0] r4575_out;
	wire [31:0] r4576_out;
	wire [31:0] r4577_out;
	wire [31:0] r4578_out;
	wire [31:0] r4579_out;
	wire [31:0] r4580_out;
	wire [31:0] r4581_out;
	wire [31:0] r4582_out;
	wire [31:0] r4583_out;
	wire [31:0] r4584_out;
	wire [31:0] r4585_out;
	wire [31:0] r4586_out;
	wire [31:0] r4587_out;
	wire [31:0] r4588_out;
	wire [31:0] r4589_out;
	wire [31:0] r4590_out;
	wire [31:0] r4591_out;
	wire [31:0] r4592_out;
	wire [31:0] r4593_out;
	wire [31:0] r4594_out;
	wire [31:0] r4595_out;
	wire [31:0] r4596_out;
	wire [31:0] r4597_out;
	wire [31:0] r4598_out;
	wire [31:0] r4599_out;
	wire [31:0] r4600_out;
	wire [31:0] r4601_out;
	wire [31:0] r4602_out;
	wire [31:0] r4603_out;
	wire [31:0] r4604_out;
	wire [31:0] r4605_out;
	wire [31:0] r4606_out;
	wire [31:0] r4607_out;
	wire [31:0] r4608_out;
	wire [31:0] r4609_out;
	wire [31:0] r4610_out;
	wire [31:0] r4611_out;
	wire [31:0] r4612_out;
	wire [31:0] r4613_out;
	wire [31:0] r4614_out;
	wire [31:0] r4615_out;
	wire [31:0] r4616_out;
	wire [31:0] r4617_out;
	wire [31:0] r4618_out;
	wire [31:0] r4619_out;
	wire [31:0] r4620_out;
	wire [31:0] r4621_out;
	wire [31:0] r4622_out;
	wire [31:0] r4623_out;
	wire [31:0] r4624_out;
	wire [31:0] r4625_out;
	wire [31:0] r4626_out;
	wire [31:0] r4627_out;
	wire [31:0] r4628_out;
	wire [31:0] r4629_out;
	wire [31:0] r4630_out;
	wire [31:0] r4631_out;
	wire [31:0] r4632_out;
	wire [31:0] r4633_out;
	wire [31:0] r4634_out;
	wire [31:0] r4635_out;
	wire [31:0] r4636_out;
	wire [31:0] r4637_out;
	wire [31:0] r4638_out;
	wire [31:0] r4639_out;
	wire [31:0] r4640_out;
	wire [31:0] r4641_out;
	wire [31:0] r4642_out;
	wire [31:0] r4643_out;
	wire [31:0] r4644_out;
	wire [31:0] r4645_out;
	wire [31:0] r4646_out;
	wire [31:0] r4647_out;
	wire [31:0] r4648_out;
	wire [31:0] r4649_out;
	wire [31:0] r4650_out;
	wire [31:0] r4651_out;
	wire [31:0] r4652_out;
	wire [31:0] r4653_out;
	wire [31:0] r4654_out;
	wire [31:0] r4655_out;
	wire [31:0] r4656_out;
	wire [31:0] r4657_out;
	wire [31:0] r4658_out;
	wire [31:0] r4659_out;
	wire [31:0] r4660_out;
	wire [31:0] r4661_out;
	wire [31:0] r4662_out;
	wire [31:0] r4663_out;
	wire [31:0] r4664_out;
	wire [31:0] r4665_out;
	wire [31:0] r4666_out;
	wire [31:0] r4667_out;
	wire [31:0] r4668_out;
	wire [31:0] r4669_out;
	wire [31:0] r4670_out;
	wire [31:0] r4671_out;
	wire [31:0] r4672_out;
	wire [31:0] r4673_out;
	wire [31:0] r4674_out;
	wire [31:0] r4675_out;
	wire [31:0] r4676_out;
	wire [31:0] r4677_out;
	wire [31:0] r4678_out;
	wire [31:0] r4679_out;
	wire [31:0] r4680_out;
	wire [31:0] r4681_out;
	wire [31:0] r4682_out;
	wire [31:0] r4683_out;
	wire [31:0] r4684_out;
	wire [31:0] r4685_out;
	wire [31:0] r4686_out;
	wire [31:0] r4687_out;
	wire [31:0] r4688_out;
	wire [31:0] r4689_out;
	wire [31:0] r4690_out;
	wire [31:0] r4691_out;
	wire [31:0] r4692_out;
	wire [31:0] r4693_out;
	wire [31:0] r4694_out;
	wire [31:0] r4695_out;
	wire [31:0] r4696_out;
	wire [31:0] r4697_out;
	wire [31:0] r4698_out;
	wire [31:0] r4699_out;
	wire [31:0] r4700_out;
	wire [31:0] r4701_out;
	wire [31:0] r4702_out;
	wire [31:0] r4703_out;
	wire [31:0] r4704_out;
	wire [31:0] r4705_out;
	wire [31:0] r4706_out;
	wire [31:0] r4707_out;
	wire [31:0] r4708_out;
	wire [31:0] r4709_out;
	wire [31:0] r4710_out;
	wire [31:0] r4711_out;
	wire [31:0] r4712_out;
	wire [31:0] r4713_out;
	wire [31:0] r4714_out;
	wire [31:0] r4715_out;
	wire [31:0] r4716_out;
	wire [31:0] r4717_out;
	wire [31:0] r4718_out;
	wire [31:0] r4719_out;
	wire [31:0] r4720_out;
	wire [31:0] r4721_out;
	wire [31:0] r4722_out;
	wire [31:0] r4723_out;
	wire [31:0] r4724_out;
	wire [31:0] r4725_out;
	wire [31:0] r4726_out;
	wire [31:0] r4727_out;
	wire [31:0] r4728_out;
	wire [31:0] r4729_out;
	wire [31:0] r4730_out;
	wire [31:0] r4731_out;
	wire [31:0] r4732_out;
	wire [31:0] r4733_out;
	wire [31:0] r4734_out;
	wire [31:0] r4735_out;
	wire [31:0] r4736_out;
	wire [31:0] r4737_out;
	wire [31:0] r4738_out;
	wire [31:0] r4739_out;
	wire [31:0] r4740_out;
	wire [31:0] r4741_out;
	wire [31:0] r4742_out;
	wire [31:0] r4743_out;
	wire [31:0] r4744_out;
	wire [31:0] r4745_out;
	wire [31:0] r4746_out;
	wire [31:0] r4747_out;
	wire [31:0] r4748_out;
	wire [31:0] r4749_out;
	wire [31:0] r4750_out;
	wire [31:0] r4751_out;
	wire [31:0] r4752_out;
	wire [31:0] r4753_out;
	wire [31:0] r4754_out;
	wire [31:0] r4755_out;
	wire [31:0] r4756_out;
	wire [31:0] r4757_out;
	wire [31:0] r4758_out;
	wire [31:0] r4759_out;
	wire [31:0] r4760_out;
	wire [31:0] r4761_out;
	wire [31:0] r4762_out;
	wire [31:0] r4763_out;
	wire [31:0] r4764_out;
	wire [31:0] r4765_out;
	wire [31:0] r4766_out;
	wire [31:0] r4767_out;
	wire [31:0] r4768_out;
	wire [31:0] r4769_out;
	wire [31:0] r4770_out;
	wire [31:0] r4771_out;
	wire [31:0] r4772_out;
	wire [31:0] r4773_out;
	wire [31:0] r4774_out;
	wire [31:0] r4775_out;
	wire [31:0] r4776_out;
	wire [31:0] r4777_out;
	wire [31:0] r4778_out;
	wire [31:0] r4779_out;
	wire [31:0] r4780_out;
	wire [31:0] r4781_out;
	wire [31:0] r4782_out;
	wire [31:0] r4783_out;
	wire [31:0] r4784_out;
	wire [31:0] r4785_out;
	wire [31:0] r4786_out;
	wire [31:0] r4787_out;
	wire [31:0] r4788_out;
	wire [31:0] r4789_out;
	wire [31:0] r4790_out;
	wire [31:0] r4791_out;
	wire [31:0] r4792_out;
	wire [31:0] r4793_out;
	wire [31:0] r4794_out;
	wire [31:0] r4795_out;
	wire [31:0] r4796_out;
	wire [31:0] r4797_out;
	wire [31:0] r4798_out;
	wire [31:0] r4799_out;
	wire [31:0] r4800_out;
	wire [31:0] r4801_out;
	wire [31:0] r4802_out;
	wire [31:0] r4803_out;
	wire [31:0] r4804_out;
	wire [31:0] r4805_out;
	wire [31:0] r4806_out;
	wire [31:0] r4807_out;
	wire [31:0] r4808_out;
	wire [31:0] r4809_out;
	wire [31:0] r4810_out;
	wire [31:0] r4811_out;
	wire [31:0] r4812_out;
	wire [31:0] r4813_out;
	wire [31:0] r4814_out;
	wire [31:0] r4815_out;
	wire [31:0] r4816_out;
	wire [31:0] r4817_out;
	wire [31:0] r4818_out;
	wire [31:0] r4819_out;
	wire [31:0] r4820_out;
	wire [31:0] r4821_out;
	wire [31:0] r4822_out;
	wire [31:0] r4823_out;
	wire [31:0] r4824_out;
	wire [31:0] r4825_out;
	wire [31:0] r4826_out;
	wire [31:0] r4827_out;
	wire [31:0] r4828_out;
	wire [31:0] r4829_out;
	wire [31:0] r4830_out;
	wire [31:0] r4831_out;
	wire [31:0] r4832_out;
	wire [31:0] r4833_out;
	wire [31:0] r4834_out;
	wire [31:0] r4835_out;
	wire [31:0] r4836_out;
	wire [31:0] r4837_out;
	wire [31:0] r4838_out;
	wire [31:0] r4839_out;
	wire [31:0] r4840_out;
	wire [31:0] r4841_out;
	wire [31:0] r4842_out;
	wire [31:0] r4843_out;
	wire [31:0] r4844_out;
	wire [31:0] r4845_out;
	wire [31:0] r4846_out;
	wire [31:0] r4847_out;
	wire [31:0] r4848_out;
	wire [31:0] r4849_out;
	wire [31:0] r4850_out;
	wire [31:0] r4851_out;
	wire [31:0] r4852_out;
	wire [31:0] r4853_out;
	wire [31:0] r4854_out;
	wire [31:0] r4855_out;
	wire [31:0] r4856_out;
	wire [31:0] r4857_out;
	wire [31:0] r4858_out;
	wire [31:0] r4859_out;
	wire [31:0] r4860_out;
	wire [31:0] r4861_out;
	wire [31:0] r4862_out;
	wire [31:0] r4863_out;
	wire [31:0] r4864_out;
	wire [31:0] r4865_out;
	wire [31:0] r4866_out;
	wire [31:0] r4867_out;
	wire [31:0] r4868_out;
	wire [31:0] r4869_out;
	wire [31:0] r4870_out;
	wire [31:0] r4871_out;
	wire [31:0] r4872_out;
	wire [31:0] r4873_out;
	wire [31:0] r4874_out;
	wire [31:0] r4875_out;
	wire [31:0] r4876_out;
	wire [31:0] r4877_out;
	wire [31:0] r4878_out;
	wire [31:0] r4879_out;
	wire [31:0] r4880_out;
	wire [31:0] r4881_out;
	wire [31:0] r4882_out;
	wire [31:0] r4883_out;
	wire [31:0] r4884_out;
	wire [31:0] r4885_out;
	wire [31:0] r4886_out;
	wire [31:0] r4887_out;
	wire [31:0] r4888_out;
	wire [31:0] r4889_out;
	wire [31:0] r4890_out;
	wire [31:0] r4891_out;
	wire [31:0] r4892_out;
	wire [31:0] r4893_out;
	wire [31:0] r4894_out;
	wire [31:0] r4895_out;
	wire [31:0] r4896_out;
	wire [31:0] r4897_out;
	wire [31:0] r4898_out;
	wire [31:0] r4899_out;
	wire [31:0] r4900_out;
	wire [31:0] r4901_out;
	wire [31:0] r4902_out;
	wire [31:0] r4903_out;
	wire [31:0] r4904_out;
	wire [31:0] r4905_out;
	wire [31:0] r4906_out;
	wire [31:0] r4907_out;
	wire [31:0] r4908_out;
	wire [31:0] r4909_out;
	wire [31:0] r4910_out;
	wire [31:0] r4911_out;
	wire [31:0] r4912_out;
	wire [31:0] r4913_out;
	wire [31:0] r4914_out;
	wire [31:0] r4915_out;
	wire [31:0] r4916_out;
	wire [31:0] r4917_out;
	wire [31:0] r4918_out;
	wire [31:0] r4919_out;
	wire [31:0] r4920_out;
	wire [31:0] r4921_out;
	wire [31:0] r4922_out;
	wire [31:0] r4923_out;
	wire [31:0] r4924_out;
	wire [31:0] r4925_out;
	wire [31:0] r4926_out;
	wire [31:0] r4927_out;
	wire [31:0] r4928_out;
	wire [31:0] r4929_out;
	wire [31:0] r4930_out;
	wire [31:0] r4931_out;
	wire [31:0] r4932_out;
	wire [31:0] r4933_out;
	wire [31:0] r4934_out;
	wire [31:0] r4935_out;
	wire [31:0] r4936_out;
	wire [31:0] r4937_out;
	wire [31:0] r4938_out;
	wire [31:0] r4939_out;
	wire [31:0] r4940_out;
	wire [31:0] r4941_out;
	wire [31:0] r4942_out;
	wire [31:0] r4943_out;
	wire [31:0] r4944_out;
	wire [31:0] r4945_out;
	wire [31:0] r4946_out;
	wire [31:0] r4947_out;
	wire [31:0] r4948_out;
	wire [31:0] r4949_out;
	wire [31:0] r4950_out;
	wire [31:0] r4951_out;
	wire [31:0] r4952_out;
	wire [31:0] r4953_out;
	wire [31:0] r4954_out;
	wire [31:0] r4955_out;
	wire [31:0] r4956_out;
	wire [31:0] r4957_out;
	wire [31:0] r4958_out;
	wire [31:0] r4959_out;
	wire [31:0] r4960_out;
	wire [31:0] r4961_out;
	wire [31:0] r4962_out;
	wire [31:0] r4963_out;
	wire [31:0] r4964_out;
	wire [31:0] r4965_out;
	wire [31:0] r4966_out;
	wire [31:0] r4967_out;
	wire [31:0] r4968_out;
	wire [31:0] r4969_out;
	wire [31:0] r4970_out;
	wire [31:0] r4971_out;
	wire [31:0] r4972_out;
	wire [31:0] r4973_out;
	wire [31:0] r4974_out;
	wire [31:0] r4975_out;
	wire [31:0] r4976_out;
	wire [31:0] r4977_out;
	wire [31:0] r4978_out;
	wire [31:0] r4979_out;
	wire [31:0] r4980_out;
	wire [31:0] r4981_out;
	wire [31:0] r4982_out;
	wire [31:0] r4983_out;
	wire [31:0] r4984_out;
	wire [31:0] r4985_out;
	wire [31:0] r4986_out;
	wire [31:0] r4987_out;
	wire [31:0] r4988_out;
	wire [31:0] r4989_out;
	wire [31:0] r4990_out;
	wire [31:0] r4991_out;
	wire [31:0] r4992_out;
	wire [31:0] r4993_out;
	wire [31:0] r4994_out;
	wire [31:0] r4995_out;
	wire [31:0] r4996_out;
	wire [31:0] r4997_out;
	wire [31:0] r4998_out;
	wire [31:0] r4999_out;
	wire [31:0] r5000_out;
	wire [31:0] r5001_out;
	wire [31:0] r5002_out;
	wire [31:0] r5003_out;
	wire [31:0] r5004_out;
	wire [31:0] r5005_out;
	wire [31:0] r5006_out;
	wire [31:0] r5007_out;
	wire [31:0] r5008_out;
	wire [31:0] r5009_out;
	wire [31:0] r5010_out;
	wire [31:0] r5011_out;
	wire [31:0] r5012_out;
	wire [31:0] r5013_out;
	wire [31:0] r5014_out;
	wire [31:0] r5015_out;
	wire [31:0] r5016_out;
	wire [31:0] r5017_out;
	wire [31:0] r5018_out;
	wire [31:0] r5019_out;
	wire [31:0] r5020_out;
	wire [31:0] r5021_out;
	wire [31:0] r5022_out;
	wire [31:0] r5023_out;
	wire [31:0] r5024_out;
	wire [31:0] r5025_out;
	wire [31:0] r5026_out;
	wire [31:0] r5027_out;
	wire [31:0] r5028_out;
	wire [31:0] r5029_out;
	wire [31:0] r5030_out;
	wire [31:0] r5031_out;
	wire [31:0] r5032_out;
	wire [31:0] r5033_out;
	wire [31:0] r5034_out;
	wire [31:0] r5035_out;
	wire [31:0] r5036_out;
	wire [31:0] r5037_out;
	wire [31:0] r5038_out;
	wire [31:0] r5039_out;
	wire [31:0] r5040_out;
	wire [31:0] r5041_out;
	wire [31:0] r5042_out;
	wire [31:0] r5043_out;
	wire [31:0] r5044_out;
	wire [31:0] r5045_out;
	wire [31:0] r5046_out;
	wire [31:0] r5047_out;
	wire [31:0] r5048_out;
	wire [31:0] r5049_out;
	wire [31:0] r5050_out;
	wire [31:0] r5051_out;
	wire [31:0] r5052_out;
	wire [31:0] r5053_out;
	wire [31:0] r5054_out;
	wire [31:0] r5055_out;
	wire [31:0] r5056_out;
	wire [31:0] r5057_out;
	wire [31:0] r5058_out;
	wire [31:0] r5059_out;
	wire [31:0] r5060_out;
	wire [31:0] r5061_out;
	wire [31:0] r5062_out;
	wire [31:0] r5063_out;
	wire [31:0] r5064_out;
	wire [31:0] r5065_out;
	wire [31:0] r5066_out;
	wire [31:0] r5067_out;
	wire [31:0] r5068_out;
	wire [31:0] r5069_out;
	wire [31:0] r5070_out;
	wire [31:0] r5071_out;
	wire [31:0] r5072_out;
	wire [31:0] r5073_out;
	wire [31:0] r5074_out;
	wire [31:0] r5075_out;
	wire [31:0] r5076_out;
	wire [31:0] r5077_out;
	wire [31:0] r5078_out;
	wire [31:0] r5079_out;
	wire [31:0] r5080_out;
	wire [31:0] r5081_out;
	wire [31:0] r5082_out;
	wire [31:0] r5083_out;
	wire [31:0] r5084_out;
	wire [31:0] r5085_out;
	wire [31:0] r5086_out;
	wire [31:0] r5087_out;
	wire [31:0] r5088_out;
	wire [31:0] r5089_out;
	wire [31:0] r5090_out;
	wire [31:0] r5091_out;
	wire [31:0] r5092_out;
	wire [31:0] r5093_out;
	wire [31:0] r5094_out;
	wire [31:0] r5095_out;
	wire [31:0] r5096_out;
	wire [31:0] r5097_out;
	wire [31:0] r5098_out;
	wire [31:0] r5099_out;
	wire [31:0] r5100_out;
	wire [31:0] r5101_out;
	wire [31:0] r5102_out;
	wire [31:0] r5103_out;
	wire [31:0] r5104_out;
	wire [31:0] r5105_out;
	wire [31:0] r5106_out;
	wire [31:0] r5107_out;
	wire [31:0] r5108_out;
	wire [31:0] r5109_out;
	wire [31:0] r5110_out;
	wire [31:0] r5111_out;
	wire [31:0] r5112_out;
	wire [31:0] r5113_out;
	wire [31:0] r5114_out;
	wire [31:0] r5115_out;
	wire [31:0] r5116_out;
	wire [31:0] r5117_out;
	wire [31:0] r5118_out;
	wire [31:0] r5119_out;
	wire [31:0] r5120_out;
	wire [31:0] r5121_out;
	wire [31:0] r5122_out;
	wire [31:0] r5123_out;
	wire [31:0] r5124_out;
	wire [31:0] r5125_out;
	wire [31:0] r5126_out;
	wire [31:0] r5127_out;
	wire [31:0] r5128_out;
	wire [31:0] r5129_out;
	wire [31:0] r5130_out;
	wire [31:0] r5131_out;
	wire [31:0] r5132_out;
	wire [31:0] r5133_out;
	wire [31:0] r5134_out;
	wire [31:0] r5135_out;
	wire [31:0] r5136_out;
	wire [31:0] r5137_out;
	wire [31:0] r5138_out;
	wire [31:0] r5139_out;
	wire [31:0] r5140_out;
	wire [31:0] r5141_out;
	wire [31:0] r5142_out;
	wire [31:0] r5143_out;
	wire [31:0] r5144_out;
	wire [31:0] r5145_out;
	wire [31:0] r5146_out;
	wire [31:0] r5147_out;
	wire [31:0] r5148_out;
	wire [31:0] r5149_out;
	wire [31:0] r5150_out;
	wire [31:0] r5151_out;
	wire [31:0] r5152_out;
	wire [31:0] r5153_out;
	wire [31:0] r5154_out;
	wire [31:0] r5155_out;
	wire [31:0] r5156_out;
	wire [31:0] r5157_out;
	wire [31:0] r5158_out;
	wire [31:0] r5159_out;
	wire [31:0] r5160_out;
	wire [31:0] r5161_out;
	wire [31:0] r5162_out;
	wire [31:0] r5163_out;
	wire [31:0] r5164_out;
	wire [31:0] r5165_out;
	wire [31:0] r5166_out;
	wire [31:0] r5167_out;
	wire [31:0] r5168_out;
	wire [31:0] r5169_out;
	wire [31:0] r5170_out;
	wire [31:0] r5171_out;
	wire [31:0] r5172_out;
	wire [31:0] r5173_out;
	wire [31:0] r5174_out;
	wire [31:0] r5175_out;
	wire [31:0] r5176_out;
	wire [31:0] r5177_out;
	wire [31:0] r5178_out;
	wire [31:0] r5179_out;
	wire [31:0] r5180_out;
	wire [31:0] r5181_out;
	wire [31:0] r5182_out;
	wire [31:0] r5183_out;
	wire [31:0] r5184_out;
	wire [31:0] r5185_out;
	wire [31:0] r5186_out;
	wire [31:0] r5187_out;
	wire [31:0] r5188_out;
	wire [31:0] r5189_out;
	wire [31:0] r5190_out;
	wire [31:0] r5191_out;
	wire [31:0] r5192_out;
	wire [31:0] r5193_out;
	wire [31:0] r5194_out;
	wire [31:0] r5195_out;
	wire [31:0] r5196_out;
	wire [31:0] r5197_out;
	wire [31:0] r5198_out;
	wire [31:0] r5199_out;
	wire [31:0] r5200_out;
	wire [31:0] r5201_out;
	wire [31:0] r5202_out;
	wire [31:0] r5203_out;
	wire [31:0] r5204_out;
	wire [31:0] r5205_out;
	wire [31:0] r5206_out;
	wire [31:0] r5207_out;
	wire [31:0] r5208_out;
	wire [31:0] r5209_out;
	wire [31:0] r5210_out;
	wire [31:0] r5211_out;
	wire [31:0] r5212_out;
	wire [31:0] r5213_out;
	wire [31:0] r5214_out;
	wire [31:0] r5215_out;
	wire [31:0] r5216_out;
	wire [31:0] r5217_out;
	wire [31:0] r5218_out;
	wire [31:0] r5219_out;
	wire [31:0] r5220_out;
	wire [31:0] r5221_out;
	wire [31:0] r5222_out;
	wire [31:0] r5223_out;
	wire [31:0] r5224_out;
	wire [31:0] r5225_out;
	wire [31:0] r5226_out;
	wire [31:0] r5227_out;
	wire [31:0] r5228_out;
	wire [31:0] r5229_out;
	wire [31:0] r5230_out;
	wire [31:0] r5231_out;
	wire [31:0] r5232_out;
	wire [31:0] r5233_out;
	wire [31:0] r5234_out;
	wire [31:0] r5235_out;
	wire [31:0] r5236_out;
	wire [31:0] r5237_out;
	wire [31:0] r5238_out;
	wire [31:0] r5239_out;
	wire [31:0] r5240_out;
	wire [31:0] r5241_out;
	wire [31:0] r5242_out;
	wire [31:0] r5243_out;
	wire [31:0] r5244_out;
	wire [31:0] r5245_out;
	wire [31:0] r5246_out;
	wire [31:0] r5247_out;
	wire [31:0] r5248_out;
	wire [31:0] r5249_out;
	wire [31:0] r5250_out;
	wire [31:0] r5251_out;
	wire [31:0] r5252_out;
	wire [31:0] r5253_out;
	wire [31:0] r5254_out;
	wire [31:0] r5255_out;
	wire [31:0] r5256_out;
	wire [31:0] r5257_out;
	wire [31:0] r5258_out;
	wire [31:0] r5259_out;
	wire [31:0] r5260_out;
	wire [31:0] r5261_out;
	wire [31:0] r5262_out;
	wire [31:0] r5263_out;
	wire [31:0] r5264_out;
	wire [31:0] r5265_out;
	wire [31:0] r5266_out;
	wire [31:0] r5267_out;
	wire [31:0] r5268_out;
	wire [31:0] r5269_out;
	wire [31:0] r5270_out;
	wire [31:0] r5271_out;
	wire [31:0] r5272_out;
	wire [31:0] r5273_out;
	wire [31:0] r5274_out;
	wire [31:0] r5275_out;
	wire [31:0] r5276_out;
	wire [31:0] r5277_out;
	wire [31:0] r5278_out;
	wire [31:0] r5279_out;
	wire [31:0] r5280_out;
	wire [31:0] r5281_out;
	wire [31:0] r5282_out;
	wire [31:0] r5283_out;
	wire [31:0] r5284_out;
	wire [31:0] r5285_out;
	wire [31:0] r5286_out;
	wire [31:0] r5287_out;
	wire [31:0] r5288_out;
	wire [31:0] r5289_out;
	wire [31:0] r5290_out;
	wire [31:0] r5291_out;
	wire [31:0] r5292_out;
	wire [31:0] r5293_out;
	wire [31:0] r5294_out;
	wire [31:0] r5295_out;
	wire [31:0] r5296_out;
	wire [31:0] r5297_out;
	wire [31:0] r5298_out;
	wire [31:0] r5299_out;
	wire [31:0] r5300_out;
	wire [31:0] r5301_out;
	wire [31:0] r5302_out;
	wire [31:0] r5303_out;
	wire [31:0] r5304_out;
	wire [31:0] r5305_out;
	wire [31:0] r5306_out;
	wire [31:0] r5307_out;
	wire [31:0] r5308_out;
	wire [31:0] r5309_out;
	wire [31:0] r5310_out;
	wire [31:0] r5311_out;
	wire [31:0] r5312_out;
	wire [31:0] r5313_out;
	wire [31:0] r5314_out;
	wire [31:0] r5315_out;
	wire [31:0] r5316_out;
	wire [31:0] r5317_out;
	wire [31:0] r5318_out;
	wire [31:0] r5319_out;
	wire [31:0] r5320_out;
	wire [31:0] r5321_out;
	wire [31:0] r5322_out;
	wire [31:0] r5323_out;
	wire [31:0] r5324_out;
	wire [31:0] r5325_out;
	wire [31:0] r5326_out;
	wire [31:0] r5327_out;
	wire [31:0] r5328_out;
	wire [31:0] r5329_out;
	wire [31:0] r5330_out;
	wire [31:0] r5331_out;
	wire [31:0] r5332_out;
	wire [31:0] r5333_out;
	wire [31:0] r5334_out;
	wire [31:0] r5335_out;
	wire [31:0] r5336_out;
	wire [31:0] r5337_out;
	wire [31:0] r5338_out;
	wire [31:0] r5339_out;
	wire [31:0] r5340_out;
	wire [31:0] r5341_out;
	wire [31:0] r5342_out;
	wire [31:0] r5343_out;
	wire [31:0] r5344_out;
	wire [31:0] r5345_out;
	wire [31:0] r5346_out;
	wire [31:0] r5347_out;
	wire [31:0] r5348_out;
	wire [31:0] r5349_out;
	wire [31:0] r5350_out;
	wire [31:0] r5351_out;
	wire [31:0] r5352_out;
	wire [31:0] r5353_out;
	wire [31:0] r5354_out;
	wire [31:0] r5355_out;
	wire [31:0] r5356_out;
	wire [31:0] r5357_out;
	wire [31:0] r5358_out;
	wire [31:0] r5359_out;
	wire [31:0] r5360_out;
	wire [31:0] r5361_out;
	wire [31:0] r5362_out;
	wire [31:0] r5363_out;
	wire [31:0] r5364_out;
	wire [31:0] r5365_out;
	wire [31:0] r5366_out;
	wire [31:0] r5367_out;
	wire [31:0] r5368_out;
	wire [31:0] r5369_out;
	wire [31:0] r5370_out;
	wire [31:0] r5371_out;
	wire [31:0] r5372_out;
	wire [31:0] r5373_out;
	wire [31:0] r5374_out;
	wire [31:0] r5375_out;
	wire [31:0] r5376_out;
	wire [31:0] r5377_out;
	wire [31:0] r5378_out;
	wire [31:0] r5379_out;
	wire [31:0] r5380_out;
	wire [31:0] r5381_out;
	wire [31:0] r5382_out;
	wire [31:0] r5383_out;
	wire [31:0] r5384_out;
	wire [31:0] r5385_out;
	wire [31:0] r5386_out;
	wire [31:0] r5387_out;
	wire [31:0] r5388_out;
	wire [31:0] r5389_out;
	wire [31:0] r5390_out;
	wire [31:0] r5391_out;
	wire [31:0] r5392_out;
	wire [31:0] r5393_out;
	wire [31:0] r5394_out;
	wire [31:0] r5395_out;
	wire [31:0] r5396_out;
	wire [31:0] r5397_out;
	wire [31:0] r5398_out;
	wire [31:0] r5399_out;
	wire [31:0] r5400_out;
	wire [31:0] r5401_out;
	wire [31:0] r5402_out;
	wire [31:0] r5403_out;
	wire [31:0] r5404_out;
	wire [31:0] r5405_out;
	wire [31:0] r5406_out;
	wire [31:0] r5407_out;
	wire [31:0] r5408_out;
	wire [31:0] r5409_out;
	wire [31:0] r5410_out;
	wire [31:0] r5411_out;
	wire [31:0] r5412_out;
	wire [31:0] r5413_out;
	wire [31:0] r5414_out;
	wire [31:0] r5415_out;
	wire [31:0] r5416_out;
	wire [31:0] r5417_out;
	wire [31:0] r5418_out;
	wire [31:0] r5419_out;
	wire [31:0] r5420_out;
	wire [31:0] r5421_out;
	wire [31:0] r5422_out;
	wire [31:0] r5423_out;
	wire [31:0] r5424_out;
	wire [31:0] r5425_out;
	wire [31:0] r5426_out;
	wire [31:0] r5427_out;
	wire [31:0] r5428_out;
	wire [31:0] r5429_out;
	wire [31:0] r5430_out;
	wire [31:0] r5431_out;
	wire [31:0] r5432_out;
	wire [31:0] r5433_out;
	wire [31:0] r5434_out;
	wire [31:0] r5435_out;
	wire [31:0] r5436_out;
	wire [31:0] r5437_out;
	wire [31:0] r5438_out;
	wire [31:0] r5439_out;
	wire [31:0] r5440_out;
	wire [31:0] r5441_out;
	wire [31:0] r5442_out;
	wire [31:0] r5443_out;
	wire [31:0] r5444_out;
	wire [31:0] r5445_out;
	wire [31:0] r5446_out;
	wire [31:0] r5447_out;
	wire [31:0] r5448_out;
	wire [31:0] r5449_out;
	wire [31:0] r5450_out;
	wire [31:0] r5451_out;
	wire [31:0] r5452_out;
	wire [31:0] r5453_out;
	wire [31:0] r5454_out;
	wire [31:0] r5455_out;
	wire [31:0] r5456_out;
	wire [31:0] r5457_out;
	wire [31:0] r5458_out;
	wire [31:0] r5459_out;
	wire [31:0] r5460_out;
	wire [31:0] r5461_out;
	wire [31:0] r5462_out;
	wire [31:0] r5463_out;
	wire [31:0] r5464_out;
	wire [31:0] r5465_out;
	wire [31:0] r5466_out;
	wire [31:0] r5467_out;
	wire [31:0] r5468_out;
	wire [31:0] r5469_out;
	wire [31:0] r5470_out;
	wire [31:0] r5471_out;
	wire [31:0] r5472_out;
	wire [31:0] r5473_out;
	wire [31:0] r5474_out;
	wire [31:0] r5475_out;
	wire [31:0] r5476_out;
	wire [31:0] r5477_out;
	wire [31:0] r5478_out;
	wire [31:0] r5479_out;
	wire [31:0] r5480_out;
	wire [31:0] r5481_out;
	wire [31:0] r5482_out;
	wire [31:0] r5483_out;
	wire [31:0] r5484_out;
	wire [31:0] r5485_out;
	wire [31:0] r5486_out;
	wire [31:0] r5487_out;
	wire [31:0] r5488_out;
	wire [31:0] r5489_out;
	wire [31:0] r5490_out;
	wire [31:0] r5491_out;
	wire [31:0] r5492_out;
	wire [31:0] r5493_out;
	wire [31:0] r5494_out;
	wire [31:0] r5495_out;
	wire [31:0] r5496_out;
	wire [31:0] r5497_out;
	wire [31:0] r5498_out;
	wire [31:0] r5499_out;
	wire [31:0] r5500_out;
	wire [31:0] r5501_out;
	wire [31:0] r5502_out;
	wire [31:0] r5503_out;
	wire [31:0] r5504_out;
	wire [31:0] r5505_out;
	wire [31:0] r5506_out;
	wire [31:0] r5507_out;
	wire [31:0] r5508_out;
	wire [31:0] r5509_out;
	wire [31:0] r5510_out;
	wire [31:0] r5511_out;
	wire [31:0] r5512_out;
	wire [31:0] r5513_out;
	wire [31:0] r5514_out;
	wire [31:0] r5515_out;
	wire [31:0] r5516_out;
	wire [31:0] r5517_out;
	wire [31:0] r5518_out;
	wire [31:0] r5519_out;
	wire [31:0] r5520_out;
	wire [31:0] r5521_out;
	wire [31:0] r5522_out;
	wire [31:0] r5523_out;
	wire [31:0] r5524_out;
	wire [31:0] r5525_out;
	wire [31:0] r5526_out;
	wire [31:0] r5527_out;
	wire [31:0] r5528_out;
	wire [31:0] r5529_out;
	wire [31:0] r5530_out;
	wire [31:0] r5531_out;
	wire [31:0] r5532_out;
	wire [31:0] r5533_out;
	wire [31:0] r5534_out;
	wire [31:0] r5535_out;
	wire [31:0] r5536_out;
	wire [31:0] r5537_out;
	wire [31:0] r5538_out;
	wire [31:0] r5539_out;
	wire [31:0] r5540_out;
	wire [31:0] r5541_out;
	wire [31:0] r5542_out;
	wire [31:0] r5543_out;
	wire [31:0] r5544_out;
	wire [31:0] r5545_out;
	wire [31:0] r5546_out;
	wire [31:0] r5547_out;
	wire [31:0] r5548_out;
	wire [31:0] r5549_out;
	wire [31:0] r5550_out;
	wire [31:0] r5551_out;
	wire [31:0] r5552_out;
	wire [31:0] r5553_out;
	wire [31:0] r5554_out;
	wire [31:0] r5555_out;
	wire [31:0] r5556_out;
	wire [31:0] r5557_out;
	wire [31:0] r5558_out;
	wire [31:0] r5559_out;
	wire [31:0] r5560_out;
	wire [31:0] r5561_out;
	wire [31:0] r5562_out;
	wire [31:0] r5563_out;
	wire [31:0] r5564_out;
	wire [31:0] r5565_out;
	wire [31:0] r5566_out;
	wire [31:0] r5567_out;
	wire [31:0] r5568_out;
	wire [31:0] r5569_out;
	wire [31:0] r5570_out;
	wire [31:0] r5571_out;
	wire [31:0] r5572_out;
	wire [31:0] r5573_out;
	wire [31:0] r5574_out;
	wire [31:0] r5575_out;
	wire [31:0] r5576_out;
	wire [31:0] r5577_out;
	wire [31:0] r5578_out;
	wire [31:0] r5579_out;
	wire [31:0] r5580_out;
	wire [31:0] r5581_out;
	wire [31:0] r5582_out;
	wire [31:0] r5583_out;
	wire [31:0] r5584_out;
	wire [31:0] r5585_out;
	wire [31:0] r5586_out;
	wire [31:0] r5587_out;
	wire [31:0] r5588_out;
	wire [31:0] r5589_out;
	wire [31:0] r5590_out;
	wire [31:0] r5591_out;
	wire [31:0] r5592_out;
	wire [31:0] r5593_out;
	wire [31:0] r5594_out;
	wire [31:0] r5595_out;
	wire [31:0] r5596_out;
	wire [31:0] r5597_out;
	wire [31:0] r5598_out;
	wire [31:0] r5599_out;
	wire [31:0] r5600_out;
	wire [31:0] r5601_out;
	wire [31:0] r5602_out;
	wire [31:0] r5603_out;
	wire [31:0] r5604_out;
	wire [31:0] r5605_out;
	wire [31:0] r5606_out;
	wire [31:0] r5607_out;
	wire [31:0] r5608_out;
	wire [31:0] r5609_out;
	wire [31:0] r5610_out;
	wire [31:0] r5611_out;
	wire [31:0] r5612_out;
	wire [31:0] r5613_out;
	wire [31:0] r5614_out;
	wire [31:0] r5615_out;
	wire [31:0] r5616_out;
	wire [31:0] r5617_out;
	wire [31:0] r5618_out;
	wire [31:0] r5619_out;
	wire [31:0] r5620_out;
	wire [31:0] r5621_out;
	wire [31:0] r5622_out;
	wire [31:0] r5623_out;
	wire [31:0] r5624_out;
	wire [31:0] r5625_out;
	wire [31:0] r5626_out;
	wire [31:0] r5627_out;
	wire [31:0] r5628_out;
	wire [31:0] r5629_out;
	wire [31:0] r5630_out;
	wire [31:0] r5631_out;
	wire [31:0] r5632_out;
	wire [31:0] r5633_out;
	wire [31:0] r5634_out;
	wire [31:0] r5635_out;
	wire [31:0] r5636_out;
	wire [31:0] r5637_out;
	wire [31:0] r5638_out;
	wire [31:0] r5639_out;
	wire [31:0] r5640_out;
	wire [31:0] r5641_out;
	wire [31:0] r5642_out;
	wire [31:0] r5643_out;
	wire [31:0] r5644_out;
	wire [31:0] r5645_out;
	wire [31:0] r5646_out;
	wire [31:0] r5647_out;
	wire [31:0] r5648_out;
	wire [31:0] r5649_out;
	wire [31:0] r5650_out;
	wire [31:0] r5651_out;
	wire [31:0] r5652_out;
	wire [31:0] r5653_out;
	wire [31:0] r5654_out;
	wire [31:0] r5655_out;
	wire [31:0] r5656_out;
	wire [31:0] r5657_out;
	wire [31:0] r5658_out;
	wire [31:0] r5659_out;
	wire [31:0] r5660_out;
	wire [31:0] r5661_out;
	wire [31:0] r5662_out;
	wire [31:0] r5663_out;
	wire [31:0] r5664_out;
	wire [31:0] r5665_out;
	wire [31:0] r5666_out;
	wire [31:0] r5667_out;
	wire [31:0] r5668_out;
	wire [31:0] r5669_out;
	wire [31:0] r5670_out;
	wire [31:0] r5671_out;
	wire [31:0] r5672_out;
	wire [31:0] r5673_out;
	wire [31:0] r5674_out;
	wire [31:0] r5675_out;
	wire [31:0] r5676_out;
	wire [31:0] r5677_out;
	wire [31:0] r5678_out;
	wire [31:0] r5679_out;
	wire [31:0] r5680_out;
	wire [31:0] r5681_out;
	wire [31:0] r5682_out;
	wire [31:0] r5683_out;
	wire [31:0] r5684_out;
	wire [31:0] r5685_out;
	wire [31:0] r5686_out;
	wire [31:0] r5687_out;
	wire [31:0] r5688_out;
	wire [31:0] r5689_out;
	wire [31:0] r5690_out;
	wire [31:0] r5691_out;
	wire [31:0] r5692_out;
	wire [31:0] r5693_out;
	wire [31:0] r5694_out;
	wire [31:0] r5695_out;
	wire [31:0] r5696_out;
	wire [31:0] r5697_out;
	wire [31:0] r5698_out;
	wire [31:0] r5699_out;
	wire [31:0] r5700_out;
	wire [31:0] r5701_out;
	wire [31:0] r5702_out;
	wire [31:0] r5703_out;
	wire [31:0] r5704_out;
	wire [31:0] r5705_out;
	wire [31:0] r5706_out;
	wire [31:0] r5707_out;
	wire [31:0] r5708_out;
	wire [31:0] r5709_out;
	wire [31:0] r5710_out;
	wire [31:0] r5711_out;
	wire [31:0] r5712_out;
	wire [31:0] r5713_out;
	wire [31:0] r5714_out;
	wire [31:0] r5715_out;
	wire [31:0] r5716_out;
	wire [31:0] r5717_out;
	wire [31:0] r5718_out;
	wire [31:0] r5719_out;
	wire [31:0] r5720_out;
	wire [31:0] r5721_out;
	wire [31:0] r5722_out;
	wire [31:0] r5723_out;
	wire [31:0] r5724_out;
	wire [31:0] r5725_out;
	wire [31:0] r5726_out;
	wire [31:0] r5727_out;
	wire [31:0] r5728_out;
	wire [31:0] r5729_out;
	wire [31:0] r5730_out;
	wire [31:0] r5731_out;
	wire [31:0] r5732_out;
	wire [31:0] r5733_out;
	wire [31:0] r5734_out;
	wire [31:0] r5735_out;
	wire [31:0] r5736_out;
	wire [31:0] r5737_out;
	wire [31:0] r5738_out;
	wire [31:0] r5739_out;
	wire [31:0] r5740_out;
	wire [31:0] r5741_out;
	wire [31:0] r5742_out;
	wire [31:0] r5743_out;
	wire [31:0] r5744_out;
	wire [31:0] r5745_out;
	wire [31:0] r5746_out;
	wire [31:0] r5747_out;
	wire [31:0] r5748_out;
	wire [31:0] r5749_out;
	wire [31:0] r5750_out;
	wire [31:0] r5751_out;
	wire [31:0] r5752_out;
	wire [31:0] r5753_out;
	wire [31:0] r5754_out;
	wire [31:0] r5755_out;
	wire [31:0] r5756_out;
	wire [31:0] r5757_out;
	wire [31:0] r5758_out;
	wire [31:0] r5759_out;
	wire [31:0] r5760_out;
	wire [31:0] r5761_out;
	wire [31:0] r5762_out;
	wire [31:0] r5763_out;
	wire [31:0] r5764_out;
	wire [31:0] r5765_out;
	wire [31:0] r5766_out;
	wire [31:0] r5767_out;
	wire [31:0] r5768_out;
	wire [31:0] r5769_out;
	wire [31:0] r5770_out;
	wire [31:0] r5771_out;
	wire [31:0] r5772_out;
	wire [31:0] r5773_out;
	wire [31:0] r5774_out;
	wire [31:0] r5775_out;
	wire [31:0] r5776_out;
	wire [31:0] r5777_out;
	wire [31:0] r5778_out;
	wire [31:0] r5779_out;
	wire [31:0] r5780_out;
	wire [31:0] r5781_out;
	wire [31:0] r5782_out;
	wire [31:0] r5783_out;
	wire [31:0] r5784_out;
	wire [31:0] r5785_out;
	wire [31:0] r5786_out;
	wire [31:0] r5787_out;
	wire [31:0] r5788_out;
	wire [31:0] r5789_out;
	wire [31:0] r5790_out;
	wire [31:0] r5791_out;
	wire [31:0] r5792_out;
	wire [31:0] r5793_out;
	wire [31:0] r5794_out;
	wire [31:0] r5795_out;
	wire [31:0] r5796_out;
	wire [31:0] r5797_out;
	wire [31:0] r5798_out;
	wire [31:0] r5799_out;
	wire [31:0] r5800_out;
	wire [31:0] r5801_out;
	wire [31:0] r5802_out;
	wire [31:0] r5803_out;
	wire [31:0] r5804_out;
	wire [31:0] r5805_out;
	wire [31:0] r5806_out;
	wire [31:0] r5807_out;
	wire [31:0] r5808_out;
	wire [31:0] r5809_out;
	wire [31:0] r5810_out;
	wire [31:0] r5811_out;
	wire [31:0] r5812_out;
	wire [31:0] r5813_out;
	wire [31:0] r5814_out;
	wire [31:0] r5815_out;
	wire [31:0] r5816_out;
	wire [31:0] r5817_out;
	wire [31:0] r5818_out;
	wire [31:0] r5819_out;
	wire [31:0] r5820_out;
	wire [31:0] r5821_out;
	wire [31:0] r5822_out;
	wire [31:0] r5823_out;
	wire [31:0] r5824_out;
	wire [31:0] r5825_out;
	wire [31:0] r5826_out;
	wire [31:0] r5827_out;
	wire [31:0] r5828_out;
	wire [31:0] r5829_out;
	wire [31:0] r5830_out;
	wire [31:0] r5831_out;
	wire [31:0] r5832_out;
	wire [31:0] r5833_out;
	wire [31:0] r5834_out;
	wire [31:0] r5835_out;
	wire [31:0] r5836_out;
	wire [31:0] r5837_out;
	wire [31:0] r5838_out;
	wire [31:0] r5839_out;
	wire [31:0] r5840_out;
	wire [31:0] r5841_out;
	wire [31:0] r5842_out;
	wire [31:0] r5843_out;
	wire [31:0] r5844_out;
	wire [31:0] r5845_out;
	wire [31:0] r5846_out;
	wire [31:0] r5847_out;
	wire [31:0] r5848_out;
	wire [31:0] r5849_out;
	wire [31:0] r5850_out;
	wire [31:0] r5851_out;
	wire [31:0] r5852_out;
	wire [31:0] r5853_out;
	wire [31:0] r5854_out;
	wire [31:0] r5855_out;
	wire [31:0] r5856_out;
	wire [31:0] r5857_out;
	wire [31:0] r5858_out;
	wire [31:0] r5859_out;
	wire [31:0] r5860_out;
	wire [31:0] r5861_out;
	wire [31:0] r5862_out;
	wire [31:0] r5863_out;
	wire [31:0] r5864_out;
	wire [31:0] r5865_out;
	wire [31:0] r5866_out;
	wire [31:0] r5867_out;
	wire [31:0] r5868_out;
	wire [31:0] r5869_out;
	wire [31:0] r5870_out;
	wire [31:0] r5871_out;
	wire [31:0] r5872_out;
	wire [31:0] r5873_out;
	wire [31:0] r5874_out;
	wire [31:0] r5875_out;
	wire [31:0] r5876_out;
	wire [31:0] r5877_out;
	wire [31:0] r5878_out;
	wire [31:0] r5879_out;
	wire [31:0] r5880_out;
	wire [31:0] r5881_out;
	wire [31:0] r5882_out;
	wire [31:0] r5883_out;
	wire [31:0] r5884_out;
	wire [31:0] r5885_out;
	wire [31:0] r5886_out;
	wire [31:0] r5887_out;
	wire [31:0] r5888_out;
	wire [31:0] r5889_out;
	wire [31:0] r5890_out;
	wire [31:0] r5891_out;
	wire [31:0] r5892_out;
	wire [31:0] r5893_out;
	wire [31:0] r5894_out;
	wire [31:0] r5895_out;
	wire [31:0] r5896_out;
	wire [31:0] r5897_out;
	wire [31:0] r5898_out;
	wire [31:0] r5899_out;
	wire [31:0] r5900_out;
	wire [31:0] r5901_out;
	wire [31:0] r5902_out;
	wire [31:0] r5903_out;
	wire [31:0] r5904_out;
	wire [31:0] r5905_out;
	wire [31:0] r5906_out;
	wire [31:0] r5907_out;
	wire [31:0] r5908_out;
	wire [31:0] r5909_out;
	wire [31:0] r5910_out;
	wire [31:0] r5911_out;
	wire [31:0] r5912_out;
	wire [31:0] r5913_out;
	wire [31:0] r5914_out;
	wire [31:0] r5915_out;
	wire [31:0] r5916_out;
	wire [31:0] r5917_out;
	wire [31:0] r5918_out;
	wire [31:0] r5919_out;
	wire [31:0] r5920_out;
	wire [31:0] r5921_out;
	wire [31:0] r5922_out;
	wire [31:0] r5923_out;
	wire [31:0] r5924_out;
	wire [31:0] r5925_out;
	wire [31:0] r5926_out;
	wire [31:0] r5927_out;
	wire [31:0] r5928_out;
	wire [31:0] r5929_out;
	wire [31:0] r5930_out;
	wire [31:0] r5931_out;
	wire [31:0] r5932_out;
	wire [31:0] r5933_out;
	wire [31:0] r5934_out;
	wire [31:0] r5935_out;
	wire [31:0] r5936_out;
	wire [31:0] r5937_out;
	wire [31:0] r5938_out;
	wire [31:0] r5939_out;
	wire [31:0] r5940_out;
	wire [31:0] r5941_out;
	wire [31:0] r5942_out;
	wire [31:0] r5943_out;
	wire [31:0] r5944_out;
	wire [31:0] r5945_out;
	wire [31:0] r5946_out;
	wire [31:0] r5947_out;
	wire [31:0] r5948_out;
	wire [31:0] r5949_out;
	wire [31:0] r5950_out;
	wire [31:0] r5951_out;
	wire [31:0] r5952_out;
	wire [31:0] r5953_out;
	wire [31:0] r5954_out;
	wire [31:0] r5955_out;
	wire [31:0] r5956_out;
	wire [31:0] r5957_out;
	wire [31:0] r5958_out;
	wire [31:0] r5959_out;
	wire [31:0] r5960_out;
	wire [31:0] r5961_out;
	wire [31:0] r5962_out;
	wire [31:0] r5963_out;
	wire [31:0] r5964_out;
	wire [31:0] r5965_out;
	wire [31:0] r5966_out;
	wire [31:0] r5967_out;
	wire [31:0] r5968_out;
	wire [31:0] r5969_out;
	wire [31:0] r5970_out;
	wire [31:0] r5971_out;
	wire [31:0] r5972_out;
	wire [31:0] r5973_out;
	wire [31:0] r5974_out;
	wire [31:0] r5975_out;
	wire [31:0] r5976_out;
	wire [31:0] r5977_out;
	wire [31:0] r5978_out;
	wire [31:0] r5979_out;
	wire [31:0] r5980_out;
	wire [31:0] r5981_out;
	wire [31:0] r5982_out;
	wire [31:0] r5983_out;
	wire [31:0] r5984_out;
	wire [31:0] r5985_out;
	wire [31:0] r5986_out;
	wire [31:0] r5987_out;
	wire [31:0] r5988_out;
	wire [31:0] r5989_out;
	wire [31:0] r5990_out;
	wire [31:0] r5991_out;
	wire [31:0] r5992_out;
	wire [31:0] r5993_out;
	wire [31:0] r5994_out;
	wire [31:0] r5995_out;
	wire [31:0] r5996_out;
	wire [31:0] r5997_out;
	wire [31:0] r5998_out;
	wire [31:0] r5999_out;
	wire [31:0] r6000_out;
	wire [31:0] r6001_out;
	wire [31:0] r6002_out;
	wire [31:0] r6003_out;
	wire [31:0] r6004_out;
	wire [31:0] r6005_out;
	wire [31:0] r6006_out;
	wire [31:0] r6007_out;
	wire [31:0] r6008_out;
	wire [31:0] r6009_out;
	wire [31:0] r6010_out;
	wire [31:0] r6011_out;
	wire [31:0] r6012_out;
	wire [31:0] r6013_out;
	wire [31:0] r6014_out;
	wire [31:0] r6015_out;
	wire [31:0] r6016_out;
	wire [31:0] r6017_out;
	wire [31:0] r6018_out;
	wire [31:0] r6019_out;
	wire [31:0] r6020_out;
	wire [31:0] r6021_out;
	wire [31:0] r6022_out;
	wire [31:0] r6023_out;
	wire [31:0] r6024_out;
	wire [31:0] r6025_out;
	wire [31:0] r6026_out;
	wire [31:0] r6027_out;
	wire [31:0] r6028_out;
	wire [31:0] r6029_out;
	wire [31:0] r6030_out;
	wire [31:0] r6031_out;
	wire [31:0] r6032_out;
	wire [31:0] r6033_out;
	wire [31:0] r6034_out;
	wire [31:0] r6035_out;
	wire [31:0] r6036_out;
	wire [31:0] r6037_out;
	wire [31:0] r6038_out;
	wire [31:0] r6039_out;
	wire [31:0] r6040_out;
	wire [31:0] r6041_out;
	wire [31:0] r6042_out;
	wire [31:0] r6043_out;
	wire [31:0] r6044_out;
	wire [31:0] r6045_out;
	wire [31:0] r6046_out;
	wire [31:0] r6047_out;
	wire [31:0] r6048_out;
	wire [31:0] r6049_out;
	wire [31:0] r6050_out;
	wire [31:0] r6051_out;
	wire [31:0] r6052_out;
	wire [31:0] r6053_out;
	wire [31:0] r6054_out;
	wire [31:0] r6055_out;
	wire [31:0] r6056_out;
	wire [31:0] r6057_out;
	wire [31:0] r6058_out;
	wire [31:0] r6059_out;
	wire [31:0] r6060_out;
	wire [31:0] r6061_out;
	wire [31:0] r6062_out;
	wire [31:0] r6063_out;
	wire [31:0] r6064_out;
	wire [31:0] r6065_out;
	wire [31:0] r6066_out;
	wire [31:0] r6067_out;
	wire [31:0] r6068_out;
	wire [31:0] r6069_out;
	wire [31:0] r6070_out;
	wire [31:0] r6071_out;
	wire [31:0] r6072_out;
	wire [31:0] r6073_out;
	wire [31:0] r6074_out;
	wire [31:0] r6075_out;
	wire [31:0] r6076_out;
	wire [31:0] r6077_out;
	wire [31:0] r6078_out;
	wire [31:0] r6079_out;
	wire [31:0] r6080_out;
	wire [31:0] r6081_out;
	wire [31:0] r6082_out;
	wire [31:0] r6083_out;
	wire [31:0] r6084_out;
	wire [31:0] r6085_out;
	wire [31:0] r6086_out;
	wire [31:0] r6087_out;
	wire [31:0] r6088_out;
	wire [31:0] r6089_out;
	wire [31:0] r6090_out;
	wire [31:0] r6091_out;
	wire [31:0] r6092_out;
	wire [31:0] r6093_out;
	wire [31:0] r6094_out;
	wire [31:0] r6095_out;
	wire [31:0] r6096_out;
	wire [31:0] r6097_out;
	wire [31:0] r6098_out;
	wire [31:0] r6099_out;
	wire [31:0] r6100_out;
	wire [31:0] r6101_out;
	wire [31:0] r6102_out;
	wire [31:0] r6103_out;
	wire [31:0] r6104_out;
	wire [31:0] r6105_out;
	wire [31:0] r6106_out;
	wire [31:0] r6107_out;
	wire [31:0] r6108_out;
	wire [31:0] r6109_out;
	wire [31:0] r6110_out;
	wire [31:0] r6111_out;
	wire [31:0] r6112_out;
	wire [31:0] r6113_out;
	wire [31:0] r6114_out;
	wire [31:0] r6115_out;
	wire [31:0] r6116_out;
	wire [31:0] r6117_out;
	wire [31:0] r6118_out;
	wire [31:0] r6119_out;
	wire [31:0] r6120_out;
	wire [31:0] r6121_out;
	wire [31:0] r6122_out;
	wire [31:0] r6123_out;
	wire [31:0] r6124_out;
	wire [31:0] r6125_out;
	wire [31:0] r6126_out;
	wire [31:0] r6127_out;
	wire [31:0] r6128_out;
	wire [31:0] r6129_out;
	wire [31:0] r6130_out;
	wire [31:0] r6131_out;
	wire [31:0] r6132_out;
	wire [31:0] r6133_out;
	wire [31:0] r6134_out;
	wire [31:0] r6135_out;
	wire [31:0] r6136_out;
	wire [31:0] r6137_out;
	wire [31:0] r6138_out;
	wire [31:0] r6139_out;
	wire [31:0] r6140_out;
	wire [31:0] r6141_out;
	wire [31:0] r6142_out;
	wire [31:0] r6143_out;
	wire [31:0] r6144_out;
	wire [31:0] r6145_out;
	wire [31:0] r6146_out;
	wire [31:0] r6147_out;
	wire [31:0] r6148_out;
	wire [31:0] r6149_out;
	wire [31:0] r6150_out;
	wire [31:0] r6151_out;
	wire [31:0] r6152_out;
	wire [31:0] r6153_out;
	wire [31:0] r6154_out;
	wire [31:0] r6155_out;
	wire [31:0] r6156_out;
	wire [31:0] r6157_out;
	wire [31:0] r6158_out;
	wire [31:0] r6159_out;
	wire [31:0] r6160_out;
	wire [31:0] r6161_out;
	wire [31:0] r6162_out;
	wire [31:0] r6163_out;
	wire [31:0] r6164_out;
	wire [31:0] r6165_out;
	wire [31:0] r6166_out;
	wire [31:0] r6167_out;
	wire [31:0] r6168_out;
	wire [31:0] r6169_out;
	wire [31:0] r6170_out;
	wire [31:0] r6171_out;
	wire [31:0] r6172_out;
	wire [31:0] r6173_out;
	wire [31:0] r6174_out;
	wire [31:0] r6175_out;
	wire [31:0] r6176_out;
	wire [31:0] r6177_out;
	wire [31:0] r6178_out;
	wire [31:0] r6179_out;
	wire [31:0] r6180_out;
	wire [31:0] r6181_out;
	wire [31:0] r6182_out;
	wire [31:0] r6183_out;
	wire [31:0] r6184_out;
	wire [31:0] r6185_out;
	wire [31:0] r6186_out;
	wire [31:0] r6187_out;
	wire [31:0] r6188_out;
	wire [31:0] r6189_out;
	wire [31:0] r6190_out;
	wire [31:0] r6191_out;
	wire [31:0] r6192_out;
	wire [31:0] r6193_out;
	wire [31:0] r6194_out;
	wire [31:0] r6195_out;
	wire [31:0] r6196_out;
	wire [31:0] r6197_out;
	wire [31:0] r6198_out;
	wire [31:0] r6199_out;
	wire [31:0] r6200_out;
	wire [31:0] r6201_out;
	wire [31:0] r6202_out;
	wire [31:0] r6203_out;
	wire [31:0] r6204_out;
	wire [31:0] r6205_out;
	wire [31:0] r6206_out;
	wire [31:0] r6207_out;
	wire [31:0] r6208_out;
	wire [31:0] r6209_out;
	wire [31:0] r6210_out;
	wire [31:0] r6211_out;
	wire [31:0] r6212_out;
	wire [31:0] r6213_out;
	wire [31:0] r6214_out;
	wire [31:0] r6215_out;
	wire [31:0] r6216_out;
	wire [31:0] r6217_out;
	wire [31:0] r6218_out;
	wire [31:0] r6219_out;
	wire [31:0] r6220_out;
	wire [31:0] r6221_out;
	wire [31:0] r6222_out;
	wire [31:0] r6223_out;
	wire [31:0] r6224_out;
	wire [31:0] r6225_out;
	wire [31:0] r6226_out;
	wire [31:0] r6227_out;
	wire [31:0] r6228_out;
	wire [31:0] r6229_out;
	wire [31:0] r6230_out;
	wire [31:0] r6231_out;
	wire [31:0] r6232_out;
	wire [31:0] r6233_out;
	wire [31:0] r6234_out;
	wire [31:0] r6235_out;
	wire [31:0] r6236_out;
	wire [31:0] r6237_out;
	wire [31:0] r6238_out;
	wire [31:0] r6239_out;
	wire [31:0] r6240_out;
	wire [31:0] r6241_out;
	wire [31:0] r6242_out;
	wire [31:0] r6243_out;
	wire [31:0] r6244_out;
	wire [31:0] r6245_out;
	wire [31:0] r6246_out;
	wire [31:0] r6247_out;
	wire [31:0] r6248_out;
	wire [31:0] r6249_out;
	wire [31:0] r6250_out;
	wire [31:0] r6251_out;
	wire [31:0] r6252_out;
	wire [31:0] r6253_out;
	wire [31:0] r6254_out;
	wire [31:0] r6255_out;
	wire [31:0] r6256_out;
	wire [31:0] r6257_out;
	wire [31:0] r6258_out;
	wire [31:0] r6259_out;
	wire [31:0] r6260_out;
	wire [31:0] r6261_out;
	wire [31:0] r6262_out;
	wire [31:0] r6263_out;
	wire [31:0] r6264_out;
	wire [31:0] r6265_out;
	wire [31:0] r6266_out;
	wire [31:0] r6267_out;
	wire [31:0] r6268_out;
	wire [31:0] r6269_out;
	wire [31:0] r6270_out;
	wire [31:0] r6271_out;
	wire [31:0] r6272_out;
	wire [31:0] r6273_out;
	wire [31:0] r6274_out;
	wire [31:0] r6275_out;
	wire [31:0] r6276_out;
	wire [31:0] r6277_out;
	wire [31:0] r6278_out;
	wire [31:0] r6279_out;
	wire [31:0] r6280_out;
	wire [31:0] r6281_out;
	wire [31:0] r6282_out;
	wire [31:0] r6283_out;
	wire [31:0] r6284_out;
	wire [31:0] r6285_out;
	wire [31:0] r6286_out;
	wire [31:0] r6287_out;
	wire [31:0] r6288_out;
	wire [31:0] r6289_out;
	wire [31:0] r6290_out;
	wire [31:0] r6291_out;
	wire [31:0] r6292_out;
	wire [31:0] r6293_out;
	wire [31:0] r6294_out;
	wire [31:0] r6295_out;
	wire [31:0] r6296_out;
	wire [31:0] r6297_out;
	wire [31:0] r6298_out;
	wire [31:0] r6299_out;
	wire [31:0] r6300_out;
	wire [31:0] r6301_out;
	wire [31:0] r6302_out;
	wire [31:0] r6303_out;
	wire [31:0] r6304_out;
	wire [31:0] r6305_out;
	wire [31:0] r6306_out;
	wire [31:0] r6307_out;
	wire [31:0] r6308_out;
	wire [31:0] r6309_out;
	wire [31:0] r6310_out;
	wire [31:0] r6311_out;
	wire [31:0] r6312_out;
	wire [31:0] r6313_out;
	wire [31:0] r6314_out;
	wire [31:0] r6315_out;
	wire [31:0] r6316_out;
	wire [31:0] r6317_out;
	wire [31:0] r6318_out;
	wire [31:0] r6319_out;
	wire [31:0] r6320_out;
	wire [31:0] r6321_out;
	wire [31:0] r6322_out;
	wire [31:0] r6323_out;
	wire [31:0] r6324_out;
	wire [31:0] r6325_out;
	wire [31:0] r6326_out;
	wire [31:0] r6327_out;
	wire [31:0] r6328_out;
	wire [31:0] r6329_out;
	wire [31:0] r6330_out;
	wire [31:0] r6331_out;
	wire [31:0] r6332_out;
	wire [31:0] r6333_out;
	wire [31:0] r6334_out;
	wire [31:0] r6335_out;
	wire [31:0] r6336_out;
	wire [31:0] r6337_out;
	wire [31:0] r6338_out;
	wire [31:0] r6339_out;
	wire [31:0] r6340_out;
	wire [31:0] r6341_out;
	wire [31:0] r6342_out;
	wire [31:0] r6343_out;
	wire [31:0] r6344_out;
	wire [31:0] r6345_out;
	wire [31:0] r6346_out;
	wire [31:0] r6347_out;
	wire [31:0] r6348_out;
	wire [31:0] r6349_out;
	wire [31:0] r6350_out;
	wire [31:0] r6351_out;
	wire [31:0] r6352_out;
	wire [31:0] r6353_out;
	wire [31:0] r6354_out;
	wire [31:0] r6355_out;
	wire [31:0] r6356_out;
	wire [31:0] r6357_out;
	wire [31:0] r6358_out;
	wire [31:0] r6359_out;
	wire [31:0] r6360_out;
	wire [31:0] r6361_out;
	wire [31:0] r6362_out;
	wire [31:0] r6363_out;
	wire [31:0] r6364_out;
	wire [31:0] r6365_out;
	wire [31:0] r6366_out;
	wire [31:0] r6367_out;
	wire [31:0] r6368_out;
	wire [31:0] r6369_out;
	wire [31:0] r6370_out;
	wire [31:0] r6371_out;
	wire [31:0] r6372_out;
	wire [31:0] r6373_out;
	wire [31:0] r6374_out;
	wire [31:0] r6375_out;
	wire [31:0] r6376_out;
	wire [31:0] r6377_out;
	wire [31:0] r6378_out;
	wire [31:0] r6379_out;
	wire [31:0] r6380_out;
	wire [31:0] r6381_out;
	wire [31:0] r6382_out;
	wire [31:0] r6383_out;
	wire [31:0] r6384_out;
	wire [31:0] r6385_out;
	wire [31:0] r6386_out;
	wire [31:0] r6387_out;
	wire [31:0] r6388_out;
	wire [31:0] r6389_out;
	wire [31:0] r6390_out;
	wire [31:0] r6391_out;
	wire [31:0] r6392_out;
	wire [31:0] r6393_out;
	wire [31:0] r6394_out;
	wire [31:0] r6395_out;
	wire [31:0] r6396_out;
	wire [31:0] r6397_out;
	wire [31:0] r6398_out;
	wire [31:0] r6399_out;
	wire [31:0] r6400_out;
	wire [31:0] r6401_out;
	wire [31:0] r6402_out;
	wire [31:0] r6403_out;
	wire [31:0] r6404_out;
	wire [31:0] r6405_out;
	wire [31:0] r6406_out;
	wire [31:0] r6407_out;
	wire [31:0] r6408_out;
	wire [31:0] r6409_out;
	wire [31:0] r6410_out;
	wire [31:0] r6411_out;
	wire [31:0] r6412_out;
	wire [31:0] r6413_out;
	wire [31:0] r6414_out;
	wire [31:0] r6415_out;
	wire [31:0] r6416_out;
	wire [31:0] r6417_out;
	wire [31:0] r6418_out;
	wire [31:0] r6419_out;
	wire [31:0] r6420_out;
	wire [31:0] r6421_out;
	wire [31:0] r6422_out;
	wire [31:0] r6423_out;
	wire [31:0] r6424_out;
	wire [31:0] r6425_out;
	wire [31:0] r6426_out;
	wire [31:0] r6427_out;
	wire [31:0] r6428_out;
	wire [31:0] r6429_out;
	wire [31:0] r6430_out;
	wire [31:0] r6431_out;
	wire [31:0] r6432_out;
	wire [31:0] r6433_out;
	wire [31:0] r6434_out;
	wire [31:0] r6435_out;
	wire [31:0] r6436_out;
	wire [31:0] r6437_out;
	wire [31:0] r6438_out;
	wire [31:0] r6439_out;
	wire [31:0] r6440_out;
	wire [31:0] r6441_out;
	wire [31:0] r6442_out;
	wire [31:0] r6443_out;
	wire [31:0] r6444_out;
	wire [31:0] r6445_out;
	wire [31:0] r6446_out;
	wire [31:0] r6447_out;
	wire [31:0] r6448_out;
	wire [31:0] r6449_out;
	wire [31:0] r6450_out;
	wire [31:0] r6451_out;
	wire [31:0] r6452_out;
	wire [31:0] r6453_out;
	wire [31:0] r6454_out;
	wire [31:0] r6455_out;
	wire [31:0] r6456_out;
	wire [31:0] r6457_out;
	wire [31:0] r6458_out;
	wire [31:0] r6459_out;
	wire [31:0] r6460_out;
	wire [31:0] r6461_out;
	wire [31:0] r6462_out;
	wire [31:0] r6463_out;
	wire [31:0] r6464_out;
	wire [31:0] r6465_out;
	wire [31:0] r6466_out;
	wire [31:0] r6467_out;
	wire [31:0] r6468_out;
	wire [31:0] r6469_out;
	wire [31:0] r6470_out;
	wire [31:0] r6471_out;
	wire [31:0] r6472_out;
	wire [31:0] r6473_out;
	wire [31:0] r6474_out;
	wire [31:0] r6475_out;
	wire [31:0] r6476_out;
	wire [31:0] r6477_out;
	wire [31:0] r6478_out;
	wire [31:0] r6479_out;
	wire [31:0] r6480_out;
	wire [31:0] r6481_out;
	wire [31:0] r6482_out;
	wire [31:0] r6483_out;
	wire [31:0] r6484_out;
	wire [31:0] r6485_out;
	wire [31:0] r6486_out;
	wire [31:0] r6487_out;
	wire [31:0] r6488_out;
	wire [31:0] r6489_out;
	wire [31:0] r6490_out;
	wire [31:0] r6491_out;
	wire [31:0] r6492_out;
	wire [31:0] r6493_out;
	wire [31:0] r6494_out;
	wire [31:0] r6495_out;
	wire [31:0] r6496_out;
	wire [31:0] r6497_out;
	wire [31:0] r6498_out;
	wire [31:0] r6499_out;
	wire [31:0] r6500_out;
	wire [31:0] r6501_out;
	wire [31:0] r6502_out;
	wire [31:0] r6503_out;
	wire [31:0] r6504_out;
	wire [31:0] r6505_out;
	wire [31:0] r6506_out;
	wire [31:0] r6507_out;
	wire [31:0] r6508_out;
	wire [31:0] r6509_out;
	wire [31:0] r6510_out;
	wire [31:0] r6511_out;
	wire [31:0] r6512_out;
	wire [31:0] r6513_out;
	wire [31:0] r6514_out;
	wire [31:0] r6515_out;
	wire [31:0] r6516_out;
	wire [31:0] r6517_out;
	wire [31:0] r6518_out;
	wire [31:0] r6519_out;
	wire [31:0] r6520_out;
	wire [31:0] r6521_out;
	wire [31:0] r6522_out;
	wire [31:0] r6523_out;
	wire [31:0] r6524_out;
	wire [31:0] r6525_out;
	wire [31:0] r6526_out;
	wire [31:0] r6527_out;
	wire [31:0] r6528_out;
	wire [31:0] r6529_out;
	wire [31:0] r6530_out;
	wire [31:0] r6531_out;
	wire [31:0] r6532_out;
	wire [31:0] r6533_out;
	wire [31:0] r6534_out;
	wire [31:0] r6535_out;
	wire [31:0] r6536_out;
	wire [31:0] r6537_out;
	wire [31:0] r6538_out;
	wire [31:0] r6539_out;
	wire [31:0] r6540_out;
	wire [31:0] r6541_out;
	wire [31:0] r6542_out;
	wire [31:0] r6543_out;
	wire [31:0] r6544_out;
	wire [31:0] r6545_out;
	wire [31:0] r6546_out;
	wire [31:0] r6547_out;
	wire [31:0] r6548_out;
	wire [31:0] r6549_out;
	wire [31:0] r6550_out;
	wire [31:0] r6551_out;
	wire [31:0] r6552_out;
	wire [31:0] r6553_out;
	wire [31:0] r6554_out;
	wire [31:0] r6555_out;
	wire [31:0] r6556_out;
	wire [31:0] r6557_out;
	wire [31:0] r6558_out;
	wire [31:0] r6559_out;
	wire [31:0] r6560_out;
	wire [31:0] r6561_out;
	wire [31:0] r6562_out;
	wire [31:0] r6563_out;
	wire [31:0] r6564_out;
	wire [31:0] r6565_out;
	wire [31:0] r6566_out;
	wire [31:0] r6567_out;
	wire [31:0] r6568_out;
	wire [31:0] r6569_out;
	wire [31:0] r6570_out;
	wire [31:0] r6571_out;
	wire [31:0] r6572_out;
	wire [31:0] r6573_out;
	wire [31:0] r6574_out;
	wire [31:0] r6575_out;
	wire [31:0] r6576_out;
	wire [31:0] r6577_out;
	wire [31:0] r6578_out;
	wire [31:0] r6579_out;
	wire [31:0] r6580_out;
	wire [31:0] r6581_out;
	wire [31:0] r6582_out;
	wire [31:0] r6583_out;
	wire [31:0] r6584_out;
	wire [31:0] r6585_out;
	wire [31:0] r6586_out;
	wire [31:0] r6587_out;
	wire [31:0] r6588_out;
	wire [31:0] r6589_out;
	wire [31:0] r6590_out;
	wire [31:0] r6591_out;
	wire [31:0] r6592_out;
	wire [31:0] r6593_out;
	wire [31:0] r6594_out;
	wire [31:0] r6595_out;
	wire [31:0] r6596_out;
	wire [31:0] r6597_out;
	wire [31:0] r6598_out;
	wire [31:0] r6599_out;
	wire [31:0] r6600_out;
	wire [31:0] r6601_out;
	wire [31:0] r6602_out;
	wire [31:0] r6603_out;
	wire [31:0] r6604_out;
	wire [31:0] r6605_out;
	wire [31:0] r6606_out;
	wire [31:0] r6607_out;
	wire [31:0] r6608_out;
	wire [31:0] r6609_out;
	wire [31:0] r6610_out;
	wire [31:0] r6611_out;
	wire [31:0] r6612_out;
	wire [31:0] r6613_out;
	wire [31:0] r6614_out;
	wire [31:0] r6615_out;
	wire [31:0] r6616_out;
	wire [31:0] r6617_out;
	wire [31:0] r6618_out;
	wire [31:0] r6619_out;
	wire [31:0] r6620_out;
	wire [31:0] r6621_out;
	wire [31:0] r6622_out;
	wire [31:0] r6623_out;
	wire [31:0] r6624_out;
	wire [31:0] r6625_out;
	wire [31:0] r6626_out;
	wire [31:0] r6627_out;
	wire [31:0] r6628_out;
	wire [31:0] r6629_out;
	wire [31:0] r6630_out;
	wire [31:0] r6631_out;
	wire [31:0] r6632_out;
	wire [31:0] r6633_out;
	wire [31:0] r6634_out;
	wire [31:0] r6635_out;
	wire [31:0] r6636_out;
	wire [31:0] r6637_out;
	wire [31:0] r6638_out;
	wire [31:0] r6639_out;
	wire [31:0] r6640_out;
	wire [31:0] r6641_out;
	wire [31:0] r6642_out;
	wire [31:0] r6643_out;
	wire [31:0] r6644_out;
	wire [31:0] r6645_out;
	wire [31:0] r6646_out;
	wire [31:0] r6647_out;
	wire [31:0] r6648_out;
	wire [31:0] r6649_out;
	wire [31:0] r6650_out;
	wire [31:0] r6651_out;
	wire [31:0] r6652_out;
	wire [31:0] r6653_out;
	wire [31:0] r6654_out;
	wire [31:0] r6655_out;
	wire [31:0] r6656_out;
	wire [31:0] r6657_out;
	wire [31:0] r6658_out;
	wire [31:0] r6659_out;
	wire [31:0] r6660_out;
	wire [31:0] r6661_out;
	wire [31:0] r6662_out;
	wire [31:0] r6663_out;
	wire [31:0] r6664_out;
	wire [31:0] r6665_out;
	wire [31:0] r6666_out;
	wire [31:0] r6667_out;
	wire [31:0] r6668_out;
	wire [31:0] r6669_out;
	wire [31:0] r6670_out;
	wire [31:0] r6671_out;
	wire [31:0] r6672_out;
	wire [31:0] r6673_out;
	wire [31:0] r6674_out;
	wire [31:0] r6675_out;
	wire [31:0] r6676_out;
	wire [31:0] r6677_out;
	wire [31:0] r6678_out;
	wire [31:0] r6679_out;
	wire [31:0] r6680_out;
	wire [31:0] r6681_out;
	wire [31:0] r6682_out;
	wire [31:0] r6683_out;
	wire [31:0] r6684_out;
	wire [31:0] r6685_out;
	wire [31:0] r6686_out;
	wire [31:0] r6687_out;
	wire [31:0] r6688_out;
	wire [31:0] r6689_out;
	wire [31:0] r6690_out;
	wire [31:0] r6691_out;
	wire [31:0] r6692_out;
	wire [31:0] r6693_out;
	wire [31:0] r6694_out;
	wire [31:0] r6695_out;
	wire [31:0] r6696_out;
	wire [31:0] r6697_out;
	wire [31:0] r6698_out;
	wire [31:0] r6699_out;
	wire [31:0] r6700_out;
	wire [31:0] r6701_out;
	wire [31:0] r6702_out;
	wire [31:0] r6703_out;
	wire [31:0] r6704_out;
	wire [31:0] r6705_out;
	wire [31:0] r6706_out;
	wire [31:0] r6707_out;
	wire [31:0] r6708_out;
	wire [31:0] r6709_out;
	wire [31:0] r6710_out;
	wire [31:0] r6711_out;
	wire [31:0] r6712_out;
	wire [31:0] r6713_out;
	wire [31:0] r6714_out;
	wire [31:0] r6715_out;
	wire [31:0] r6716_out;
	wire [31:0] r6717_out;
	wire [31:0] r6718_out;
	wire [31:0] r6719_out;
	wire [31:0] r6720_out;
	wire [31:0] r6721_out;
	wire [31:0] r6722_out;
	wire [31:0] r6723_out;
	wire [31:0] r6724_out;
	wire [31:0] r6725_out;
	wire [31:0] r6726_out;
	wire [31:0] r6727_out;
	wire [31:0] r6728_out;
	wire [31:0] r6729_out;
	wire [31:0] r6730_out;
	wire [31:0] r6731_out;
	wire [31:0] r6732_out;
	wire [31:0] r6733_out;
	wire [31:0] r6734_out;
	wire [31:0] r6735_out;
	wire [31:0] r6736_out;
	wire [31:0] r6737_out;
	wire [31:0] r6738_out;
	wire [31:0] r6739_out;
	wire [31:0] r6740_out;
	wire [31:0] r6741_out;
	wire [31:0] r6742_out;
	wire [31:0] r6743_out;
	wire [31:0] r6744_out;
	wire [31:0] r6745_out;
	wire [31:0] r6746_out;
	wire [31:0] r6747_out;
	wire [31:0] r6748_out;
	wire [31:0] r6749_out;
	wire [31:0] r6750_out;
	wire [31:0] r6751_out;
	wire [31:0] r6752_out;
	wire [31:0] r6753_out;
	wire [31:0] r6754_out;
	wire [31:0] r6755_out;
	wire [31:0] r6756_out;
	wire [31:0] r6757_out;
	wire [31:0] r6758_out;
	wire [31:0] r6759_out;
	wire [31:0] r6760_out;
	wire [31:0] r6761_out;
	wire [31:0] r6762_out;
	wire [31:0] r6763_out;
	wire [31:0] r6764_out;
	wire [31:0] r6765_out;
	wire [31:0] r6766_out;
	wire [31:0] r6767_out;
	wire [31:0] r6768_out;
	wire [31:0] r6769_out;
	wire [31:0] r6770_out;
	wire [31:0] r6771_out;
	wire [31:0] r6772_out;
	wire [31:0] r6773_out;
	wire [31:0] r6774_out;
	wire [31:0] r6775_out;
	wire [31:0] r6776_out;
	wire [31:0] r6777_out;
	wire [31:0] r6778_out;
	wire [31:0] r6779_out;
	wire [31:0] r6780_out;
	wire [31:0] r6781_out;
	wire [31:0] r6782_out;
	wire [31:0] r6783_out;
	wire [31:0] r6784_out;
	wire [31:0] r6785_out;
	wire [31:0] r6786_out;
	wire [31:0] r6787_out;
	wire [31:0] r6788_out;
	wire [31:0] r6789_out;
	wire [31:0] r6790_out;
	wire [31:0] r6791_out;
	wire [31:0] r6792_out;
	wire [31:0] r6793_out;
	wire [31:0] r6794_out;
	wire [31:0] r6795_out;
	wire [31:0] r6796_out;
	wire [31:0] r6797_out;
	wire [31:0] r6798_out;
	wire [31:0] r6799_out;
	wire [31:0] r6800_out;
	wire [31:0] r6801_out;
	wire [31:0] r6802_out;
	wire [31:0] r6803_out;
	wire [31:0] r6804_out;
	wire [31:0] r6805_out;
	wire [31:0] r6806_out;
	wire [31:0] r6807_out;
	wire [31:0] r6808_out;
	wire [31:0] r6809_out;
	wire [31:0] r6810_out;
	wire [31:0] r6811_out;
	wire [31:0] r6812_out;
	wire [31:0] r6813_out;
	wire [31:0] r6814_out;
	wire [31:0] r6815_out;
	wire [31:0] r6816_out;
	wire [31:0] r6817_out;
	wire [31:0] r6818_out;
	wire [31:0] r6819_out;
	wire [31:0] r6820_out;
	wire [31:0] r6821_out;
	wire [31:0] r6822_out;
	wire [31:0] r6823_out;
	wire [31:0] r6824_out;
	wire [31:0] r6825_out;
	wire [31:0] r6826_out;
	wire [31:0] r6827_out;
	wire [31:0] r6828_out;
	wire [31:0] r6829_out;
	wire [31:0] r6830_out;
	wire [31:0] r6831_out;
	wire [31:0] r6832_out;
	wire [31:0] r6833_out;
	wire [31:0] r6834_out;
	wire [31:0] r6835_out;
	wire [31:0] r6836_out;
	wire [31:0] r6837_out;
	wire [31:0] r6838_out;
	wire [31:0] r6839_out;
	wire [31:0] r6840_out;
	wire [31:0] r6841_out;
	wire [31:0] r6842_out;
	wire [31:0] r6843_out;
	wire [31:0] r6844_out;
	wire [31:0] r6845_out;
	wire [31:0] r6846_out;
	wire [31:0] r6847_out;
	wire [31:0] r6848_out;
	wire [31:0] r6849_out;
	wire [31:0] r6850_out;
	wire [31:0] r6851_out;
	wire [31:0] r6852_out;
	wire [31:0] r6853_out;
	wire [31:0] r6854_out;
	wire [31:0] r6855_out;
	wire [31:0] r6856_out;
	wire [31:0] r6857_out;
	wire [31:0] r6858_out;
	wire [31:0] r6859_out;
	wire [31:0] r6860_out;
	wire [31:0] r6861_out;
	wire [31:0] r6862_out;
	wire [31:0] r6863_out;
	wire [31:0] r6864_out;
	wire [31:0] r6865_out;
	wire [31:0] r6866_out;
	wire [31:0] r6867_out;
	wire [31:0] r6868_out;
	wire [31:0] r6869_out;
	wire [31:0] r6870_out;
	wire [31:0] r6871_out;
	wire [31:0] r6872_out;
	wire [31:0] r6873_out;
	wire [31:0] r6874_out;
	wire [31:0] r6875_out;
	wire [31:0] r6876_out;
	wire [31:0] r6877_out;
	wire [31:0] r6878_out;
	wire [31:0] r6879_out;
	wire [31:0] r6880_out;
	wire [31:0] r6881_out;
	wire [31:0] r6882_out;
	wire [31:0] r6883_out;
	wire [31:0] r6884_out;
	wire [31:0] r6885_out;
	wire [31:0] r6886_out;
	wire [31:0] r6887_out;
	wire [31:0] r6888_out;
	wire [31:0] r6889_out;
	wire [31:0] r6890_out;
	wire [31:0] r6891_out;
	wire [31:0] r6892_out;
	wire [31:0] r6893_out;
	wire [31:0] r6894_out;
	wire [31:0] r6895_out;
	wire [31:0] r6896_out;
	wire [31:0] r6897_out;
	wire [31:0] r6898_out;
	wire [31:0] r6899_out;
	wire [31:0] r6900_out;
	wire [31:0] r6901_out;
	wire [31:0] r6902_out;
	wire [31:0] r6903_out;
	wire [31:0] r6904_out;
	wire [31:0] r6905_out;
	wire [31:0] r6906_out;
	wire [31:0] r6907_out;
	wire [31:0] r6908_out;
	wire [31:0] r6909_out;
	wire [31:0] r6910_out;
	wire [31:0] r6911_out;
	wire [31:0] r6912_out;
	wire [31:0] r6913_out;
	wire [31:0] r6914_out;
	wire [31:0] r6915_out;
	wire [31:0] r6916_out;
	wire [31:0] r6917_out;
	wire [31:0] r6918_out;
	wire [31:0] r6919_out;
	wire [31:0] r6920_out;
	wire [31:0] r6921_out;
	wire [31:0] r6922_out;
	wire [31:0] r6923_out;
	wire [31:0] r6924_out;
	wire [31:0] r6925_out;
	wire [31:0] r6926_out;
	wire [31:0] r6927_out;
	wire [31:0] r6928_out;
	wire [31:0] r6929_out;
	wire [31:0] r6930_out;
	wire [31:0] r6931_out;
	wire [31:0] r6932_out;
	wire [31:0] r6933_out;
	wire [31:0] r6934_out;
	wire [31:0] r6935_out;
	wire [31:0] r6936_out;
	wire [31:0] r6937_out;
	wire [31:0] r6938_out;
	wire [31:0] r6939_out;
	wire [31:0] r6940_out;
	wire [31:0] r6941_out;
	wire [31:0] r6942_out;
	wire [31:0] r6943_out;
	wire [31:0] r6944_out;
	wire [31:0] r6945_out;
	wire [31:0] r6946_out;
	wire [31:0] r6947_out;
	wire [31:0] r6948_out;
	wire [31:0] r6949_out;
	wire [31:0] r6950_out;
	wire [31:0] r6951_out;
	wire [31:0] r6952_out;
	wire [31:0] r6953_out;
	wire [31:0] r6954_out;
	wire [31:0] r6955_out;
	wire [31:0] r6956_out;
	wire [31:0] r6957_out;
	wire [31:0] r6958_out;
	wire [31:0] r6959_out;
	wire [31:0] r6960_out;
	wire [31:0] r6961_out;
	wire [31:0] r6962_out;
	wire [31:0] r6963_out;
	wire [31:0] r6964_out;
	wire [31:0] r6965_out;
	wire [31:0] r6966_out;
	wire [31:0] r6967_out;
	wire [31:0] r6968_out;
	wire [31:0] r6969_out;
	wire [31:0] r6970_out;
	wire [31:0] r6971_out;
	wire [31:0] r6972_out;
	wire [31:0] r6973_out;
	wire [31:0] r6974_out;
	wire [31:0] r6975_out;
	wire [31:0] r6976_out;
	wire [31:0] r6977_out;
	wire [31:0] r6978_out;
	wire [31:0] r6979_out;
	wire [31:0] r6980_out;
	wire [31:0] r6981_out;
	wire [31:0] r6982_out;
	wire [31:0] r6983_out;
	wire [31:0] r6984_out;
	wire [31:0] r6985_out;
	wire [31:0] r6986_out;
	wire [31:0] r6987_out;
	wire [31:0] r6988_out;
	wire [31:0] r6989_out;
	wire [31:0] r6990_out;
	wire [31:0] r6991_out;
	wire [31:0] r6992_out;
	wire [31:0] r6993_out;
	wire [31:0] r6994_out;
	wire [31:0] r6995_out;
	wire [31:0] r6996_out;
	wire [31:0] r6997_out;
	wire [31:0] r6998_out;
	wire [31:0] r6999_out;
	wire [31:0] r7000_out;
	wire [31:0] r7001_out;
	wire [31:0] r7002_out;
	wire [31:0] r7003_out;
	wire [31:0] r7004_out;
	wire [31:0] r7005_out;
	wire [31:0] r7006_out;
	wire [31:0] r7007_out;
	wire [31:0] r7008_out;
	wire [31:0] r7009_out;
	wire [31:0] r7010_out;
	wire [31:0] r7011_out;
	wire [31:0] r7012_out;
	wire [31:0] r7013_out;
	wire [31:0] r7014_out;
	wire [31:0] r7015_out;
	wire [31:0] r7016_out;
	wire [31:0] r7017_out;
	wire [31:0] r7018_out;
	wire [31:0] r7019_out;
	wire [31:0] r7020_out;
	wire [31:0] r7021_out;
	wire [31:0] r7022_out;
	wire [31:0] r7023_out;
	wire [31:0] r7024_out;
	wire [31:0] r7025_out;
	wire [31:0] r7026_out;
	wire [31:0] r7027_out;
	wire [31:0] r7028_out;
	wire [31:0] r7029_out;
	wire [31:0] r7030_out;
	wire [31:0] r7031_out;
	wire [31:0] r7032_out;
	wire [31:0] r7033_out;
	wire [31:0] r7034_out;
	wire [31:0] r7035_out;
	wire [31:0] r7036_out;
	wire [31:0] r7037_out;
	wire [31:0] r7038_out;
	wire [31:0] r7039_out;
	wire [31:0] r7040_out;
	wire [31:0] r7041_out;
	wire [31:0] r7042_out;
	wire [31:0] r7043_out;
	wire [31:0] r7044_out;
	wire [31:0] r7045_out;
	wire [31:0] r7046_out;
	wire [31:0] r7047_out;
	wire [31:0] r7048_out;
	wire [31:0] r7049_out;
	wire [31:0] r7050_out;
	wire [31:0] r7051_out;
	wire [31:0] r7052_out;
	wire [31:0] r7053_out;
	wire [31:0] r7054_out;
	wire [31:0] r7055_out;
	wire [31:0] r7056_out;
	wire [31:0] r7057_out;
	wire [31:0] r7058_out;
	wire [31:0] r7059_out;
	wire [31:0] r7060_out;
	wire [31:0] r7061_out;
	wire [31:0] r7062_out;
	wire [31:0] r7063_out;
	wire [31:0] r7064_out;
	wire [31:0] r7065_out;
	wire [31:0] r7066_out;
	wire [31:0] r7067_out;
	wire [31:0] r7068_out;
	wire [31:0] r7069_out;
	wire [31:0] r7070_out;
	wire [31:0] r7071_out;
	wire [31:0] r7072_out;
	wire [31:0] r7073_out;
	wire [31:0] r7074_out;
	wire [31:0] r7075_out;
	wire [31:0] r7076_out;
	wire [31:0] r7077_out;
	wire [31:0] r7078_out;
	wire [31:0] r7079_out;
	wire [31:0] r7080_out;
	wire [31:0] r7081_out;
	wire [31:0] r7082_out;
	wire [31:0] r7083_out;
	wire [31:0] r7084_out;
	wire [31:0] r7085_out;
	wire [31:0] r7086_out;
	wire [31:0] r7087_out;
	wire [31:0] r7088_out;
	wire [31:0] r7089_out;
	wire [31:0] r7090_out;
	wire [31:0] r7091_out;
	wire [31:0] r7092_out;
	wire [31:0] r7093_out;
	wire [31:0] r7094_out;
	wire [31:0] r7095_out;
	wire [31:0] r7096_out;
	wire [31:0] r7097_out;
	wire [31:0] r7098_out;
	wire [31:0] r7099_out;
	wire [31:0] r7100_out;
	wire [31:0] r7101_out;
	wire [31:0] r7102_out;
	wire [31:0] r7103_out;
	wire [31:0] r7104_out;
	wire [31:0] r7105_out;
	wire [31:0] r7106_out;
	wire [31:0] r7107_out;
	wire [31:0] r7108_out;
	wire [31:0] r7109_out;
	wire [31:0] r7110_out;
	wire [31:0] r7111_out;
	wire [31:0] r7112_out;
	wire [31:0] r7113_out;
	wire [31:0] r7114_out;
	wire [31:0] r7115_out;
	wire [31:0] r7116_out;
	wire [31:0] r7117_out;
	wire [31:0] r7118_out;
	wire [31:0] r7119_out;
	wire [31:0] r7120_out;
	wire [31:0] r7121_out;
	wire [31:0] r7122_out;
	wire [31:0] r7123_out;
	wire [31:0] r7124_out;
	wire [31:0] r7125_out;
	wire [31:0] r7126_out;
	wire [31:0] r7127_out;
	wire [31:0] r7128_out;
	wire [31:0] r7129_out;
	wire [31:0] r7130_out;
	wire [31:0] r7131_out;
	wire [31:0] r7132_out;
	wire [31:0] r7133_out;
	wire [31:0] r7134_out;
	wire [31:0] r7135_out;
	wire [31:0] r7136_out;
	wire [31:0] r7137_out;
	wire [31:0] r7138_out;
	wire [31:0] r7139_out;
	wire [31:0] r7140_out;
	wire [31:0] r7141_out;
	wire [31:0] r7142_out;
	wire [31:0] r7143_out;
	wire [31:0] r7144_out;
	wire [31:0] r7145_out;
	wire [31:0] r7146_out;
	wire [31:0] r7147_out;
	wire [31:0] r7148_out;
	wire [31:0] r7149_out;
	wire [31:0] r7150_out;
	wire [31:0] r7151_out;
	wire [31:0] r7152_out;
	wire [31:0] r7153_out;
	wire [31:0] r7154_out;
	wire [31:0] r7155_out;
	wire [31:0] r7156_out;
	wire [31:0] r7157_out;
	wire [31:0] r7158_out;
	wire [31:0] r7159_out;
	wire [31:0] r7160_out;
	wire [31:0] r7161_out;
	wire [31:0] r7162_out;
	wire [31:0] r7163_out;
	wire [31:0] r7164_out;
	wire [31:0] r7165_out;
	wire [31:0] r7166_out;
	wire [31:0] r7167_out;
	wire [31:0] r7168_out;
	wire [31:0] r7169_out;
	wire [31:0] r7170_out;
	wire [31:0] r7171_out;
	wire [31:0] r7172_out;
	wire [31:0] r7173_out;
	wire [31:0] r7174_out;
	wire [31:0] r7175_out;
	wire [31:0] r7176_out;
	wire [31:0] r7177_out;
	wire [31:0] r7178_out;
	wire [31:0] r7179_out;
	wire [31:0] r7180_out;
	wire [31:0] r7181_out;
	wire [31:0] r7182_out;
	wire [31:0] r7183_out;
	wire [31:0] r7184_out;
	wire [31:0] r7185_out;
	wire [31:0] r7186_out;
	wire [31:0] r7187_out;
	wire [31:0] r7188_out;
	wire [31:0] r7189_out;
	wire [31:0] r7190_out;
	wire [31:0] r7191_out;
	wire [31:0] r7192_out;
	wire [31:0] r7193_out;
	wire [31:0] r7194_out;
	wire [31:0] r7195_out;
	wire [31:0] r7196_out;
	wire [31:0] r7197_out;
	wire [31:0] r7198_out;
	wire [31:0] r7199_out;
	wire [31:0] r7200_out;
	wire [31:0] r7201_out;
	wire [31:0] r7202_out;
	wire [31:0] r7203_out;
	wire [31:0] r7204_out;
	wire [31:0] r7205_out;
	wire [31:0] r7206_out;
	wire [31:0] r7207_out;
	wire [31:0] r7208_out;
	wire [31:0] r7209_out;
	wire [31:0] r7210_out;
	wire [31:0] r7211_out;
	wire [31:0] r7212_out;
	wire [31:0] r7213_out;
	wire [31:0] r7214_out;
	wire [31:0] r7215_out;
	wire [31:0] r7216_out;
	wire [31:0] r7217_out;
	wire [31:0] r7218_out;
	wire [31:0] r7219_out;
	wire [31:0] r7220_out;
	wire [31:0] r7221_out;
	wire [31:0] r7222_out;
	wire [31:0] r7223_out;
	wire [31:0] r7224_out;
	wire [31:0] r7225_out;
	wire [31:0] r7226_out;
	wire [31:0] r7227_out;
	wire [31:0] r7228_out;
	wire [31:0] r7229_out;
	wire [31:0] r7230_out;
	wire [31:0] r7231_out;
	wire [31:0] r7232_out;
	wire [31:0] r7233_out;
	wire [31:0] r7234_out;
	wire [31:0] r7235_out;
	wire [31:0] r7236_out;
	wire [31:0] r7237_out;
	wire [31:0] r7238_out;
	wire [31:0] r7239_out;
	wire [31:0] r7240_out;
	wire [31:0] r7241_out;
	wire [31:0] r7242_out;
	wire [31:0] r7243_out;
	wire [31:0] r7244_out;
	wire [31:0] r7245_out;
	wire [31:0] r7246_out;
	wire [31:0] r7247_out;
	wire [31:0] r7248_out;
	wire [31:0] r7249_out;
	wire [31:0] r7250_out;
	wire [31:0] r7251_out;
	wire [31:0] r7252_out;
	wire [31:0] r7253_out;
	wire [31:0] r7254_out;
	wire [31:0] r7255_out;
	wire [31:0] r7256_out;
	wire [31:0] r7257_out;
	wire [31:0] r7258_out;
	wire [31:0] r7259_out;
	wire [31:0] r7260_out;
	wire [31:0] r7261_out;
	wire [31:0] r7262_out;
	wire [31:0] r7263_out;
	wire [31:0] r7264_out;
	wire [31:0] r7265_out;
	wire [31:0] r7266_out;
	wire [31:0] r7267_out;
	wire [31:0] r7268_out;
	wire [31:0] r7269_out;
	wire [31:0] r7270_out;
	wire [31:0] r7271_out;
	wire [31:0] r7272_out;
	wire [31:0] r7273_out;
	wire [31:0] r7274_out;
	wire [31:0] r7275_out;
	wire [31:0] r7276_out;
	wire [31:0] r7277_out;
	wire [31:0] r7278_out;
	wire [31:0] r7279_out;
	wire [31:0] r7280_out;
	wire [31:0] r7281_out;
	wire [31:0] r7282_out;
	wire [31:0] r7283_out;
	wire [31:0] r7284_out;
	wire [31:0] r7285_out;
	wire [31:0] r7286_out;
	wire [31:0] r7287_out;
	wire [31:0] r7288_out;
	wire [31:0] r7289_out;
	wire [31:0] r7290_out;
	wire [31:0] r7291_out;
	wire [31:0] r7292_out;
	wire [31:0] r7293_out;
	wire [31:0] r7294_out;
	wire [31:0] r7295_out;
	wire [31:0] r7296_out;
	wire [31:0] r7297_out;
	wire [31:0] r7298_out;
	wire [31:0] r7299_out;
	wire [31:0] r7300_out;
	wire [31:0] r7301_out;
	wire [31:0] r7302_out;
	wire [31:0] r7303_out;
	wire [31:0] r7304_out;
	wire [31:0] r7305_out;
	wire [31:0] r7306_out;
	wire [31:0] r7307_out;
	wire [31:0] r7308_out;
	wire [31:0] r7309_out;
	wire [31:0] r7310_out;
	wire [31:0] r7311_out;
	wire [31:0] r7312_out;
	wire [31:0] r7313_out;
	wire [31:0] r7314_out;
	wire [31:0] r7315_out;
	wire [31:0] r7316_out;
	wire [31:0] r7317_out;
	wire [31:0] r7318_out;
	wire [31:0] r7319_out;
	wire [31:0] r7320_out;
	wire [31:0] r7321_out;
	wire [31:0] r7322_out;
	wire [31:0] r7323_out;
	wire [31:0] r7324_out;
	wire [31:0] r7325_out;
	wire [31:0] r7326_out;
	wire [31:0] r7327_out;
	wire [31:0] r7328_out;
	wire [31:0] r7329_out;
	wire [31:0] r7330_out;
	wire [31:0] r7331_out;
	wire [31:0] r7332_out;
	wire [31:0] r7333_out;
	wire [31:0] r7334_out;
	wire [31:0] r7335_out;
	wire [31:0] r7336_out;
	wire [31:0] r7337_out;
	wire [31:0] r7338_out;
	wire [31:0] r7339_out;
	wire [31:0] r7340_out;
	wire [31:0] r7341_out;
	wire [31:0] r7342_out;
	wire [31:0] r7343_out;
	wire [31:0] r7344_out;
	wire [31:0] r7345_out;
	wire [31:0] r7346_out;
	wire [31:0] r7347_out;
	wire [31:0] r7348_out;
	wire [31:0] r7349_out;
	wire [31:0] r7350_out;
	wire [31:0] r7351_out;
	wire [31:0] r7352_out;
	wire [31:0] r7353_out;
	wire [31:0] r7354_out;
	wire [31:0] r7355_out;
	wire [31:0] r7356_out;
	wire [31:0] r7357_out;
	wire [31:0] r7358_out;
	wire [31:0] r7359_out;
	wire [31:0] r7360_out;
	wire [31:0] r7361_out;
	wire [31:0] r7362_out;
	wire [31:0] r7363_out;
	wire [31:0] r7364_out;
	wire [31:0] r7365_out;
	wire [31:0] r7366_out;
	wire [31:0] r7367_out;
	wire [31:0] r7368_out;
	wire [31:0] r7369_out;
	wire [31:0] r7370_out;
	wire [31:0] r7371_out;
	wire [31:0] r7372_out;
	wire [31:0] r7373_out;
	wire [31:0] r7374_out;
	wire [31:0] r7375_out;
	wire [31:0] r7376_out;
	wire [31:0] r7377_out;
	wire [31:0] r7378_out;
	wire [31:0] r7379_out;
	wire [31:0] r7380_out;
	wire [31:0] r7381_out;
	wire [31:0] r7382_out;
	wire [31:0] r7383_out;
	wire [31:0] r7384_out;
	wire [31:0] r7385_out;
	wire [31:0] r7386_out;
	wire [31:0] r7387_out;
	wire [31:0] r7388_out;
	wire [31:0] r7389_out;
	wire [31:0] r7390_out;
	wire [31:0] r7391_out;
	wire [31:0] r7392_out;
	wire [31:0] r7393_out;
	wire [31:0] r7394_out;
	wire [31:0] r7395_out;
	wire [31:0] r7396_out;
	wire [31:0] r7397_out;
	wire [31:0] r7398_out;
	wire [31:0] r7399_out;
	wire [31:0] r7400_out;
	wire [31:0] r7401_out;
	wire [31:0] r7402_out;
	wire [31:0] r7403_out;
	wire [31:0] r7404_out;
	wire [31:0] r7405_out;
	wire [31:0] r7406_out;
	wire [31:0] r7407_out;
	wire [31:0] r7408_out;
	wire [31:0] r7409_out;
	wire [31:0] r7410_out;
	wire [31:0] r7411_out;
	wire [31:0] r7412_out;
	wire [31:0] r7413_out;
	wire [31:0] r7414_out;
	wire [31:0] r7415_out;
	wire [31:0] r7416_out;
	wire [31:0] r7417_out;
	wire [31:0] r7418_out;
	wire [31:0] r7419_out;
	wire [31:0] r7420_out;
	wire [31:0] r7421_out;
	wire [31:0] r7422_out;
	wire [31:0] r7423_out;
	wire [31:0] r7424_out;
	wire [31:0] r7425_out;
	wire [31:0] r7426_out;
	wire [31:0] r7427_out;
	wire [31:0] r7428_out;
	wire [31:0] r7429_out;
	wire [31:0] r7430_out;
	wire [31:0] r7431_out;
	wire [31:0] r7432_out;
	wire [31:0] r7433_out;
	wire [31:0] r7434_out;
	wire [31:0] r7435_out;
	wire [31:0] r7436_out;
	wire [31:0] r7437_out;
	wire [31:0] r7438_out;
	wire [31:0] r7439_out;
	wire [31:0] r7440_out;
	wire [31:0] r7441_out;
	wire [31:0] r7442_out;
	wire [31:0] r7443_out;
	wire [31:0] r7444_out;
	wire [31:0] r7445_out;
	wire [31:0] r7446_out;
	wire [31:0] r7447_out;
	wire [31:0] r7448_out;
	wire [31:0] r7449_out;
	wire [31:0] r7450_out;
	wire [31:0] r7451_out;
	wire [31:0] r7452_out;
	wire [31:0] r7453_out;
	wire [31:0] r7454_out;
	wire [31:0] r7455_out;
	wire [31:0] r7456_out;
	wire [31:0] r7457_out;
	wire [31:0] r7458_out;
	wire [31:0] r7459_out;
	wire [31:0] r7460_out;
	wire [31:0] r7461_out;
	wire [31:0] r7462_out;
	wire [31:0] r7463_out;
	wire [31:0] r7464_out;
	wire [31:0] r7465_out;
	wire [31:0] r7466_out;
	wire [31:0] r7467_out;
	wire [31:0] r7468_out;
	wire [31:0] r7469_out;
	wire [31:0] r7470_out;
	wire [31:0] r7471_out;
	wire [31:0] r7472_out;
	wire [31:0] r7473_out;
	wire [31:0] r7474_out;
	wire [31:0] r7475_out;
	wire [31:0] r7476_out;
	wire [31:0] r7477_out;
	wire [31:0] r7478_out;
	wire [31:0] r7479_out;
	wire [31:0] r7480_out;
	wire [31:0] r7481_out;
	wire [31:0] r7482_out;
	wire [31:0] r7483_out;
	wire [31:0] r7484_out;
	wire [31:0] r7485_out;
	wire [31:0] r7486_out;
	wire [31:0] r7487_out;
	wire [31:0] r7488_out;
	wire [31:0] r7489_out;
	wire [31:0] r7490_out;
	wire [31:0] r7491_out;
	wire [31:0] r7492_out;
	wire [31:0] r7493_out;
	wire [31:0] r7494_out;
	wire [31:0] r7495_out;
	wire [31:0] r7496_out;
	wire [31:0] r7497_out;
	wire [31:0] r7498_out;
	wire [31:0] r7499_out;
	wire [31:0] r7500_out;
	wire [31:0] r7501_out;
	wire [31:0] r7502_out;
	wire [31:0] r7503_out;
	wire [31:0] r7504_out;
	wire [31:0] r7505_out;
	wire [31:0] r7506_out;
	wire [31:0] r7507_out;
	wire [31:0] r7508_out;
	wire [31:0] r7509_out;
	wire [31:0] r7510_out;
	wire [31:0] r7511_out;
	wire [31:0] r7512_out;
	wire [31:0] r7513_out;
	wire [31:0] r7514_out;
	wire [31:0] r7515_out;
	wire [31:0] r7516_out;
	wire [31:0] r7517_out;
	wire [31:0] r7518_out;
	wire [31:0] r7519_out;
	wire [31:0] r7520_out;
	wire [31:0] r7521_out;
	wire [31:0] r7522_out;
	wire [31:0] r7523_out;
	wire [31:0] r7524_out;
	wire [31:0] r7525_out;
	wire [31:0] r7526_out;
	wire [31:0] r7527_out;
	wire [31:0] r7528_out;
	wire [31:0] r7529_out;
	wire [31:0] r7530_out;
	wire [31:0] r7531_out;
	wire [31:0] r7532_out;
	wire [31:0] r7533_out;
	wire [31:0] r7534_out;
	wire [31:0] r7535_out;
	wire [31:0] r7536_out;
	wire [31:0] r7537_out;
	wire [31:0] r7538_out;
	wire [31:0] r7539_out;
	wire [31:0] r7540_out;
	wire [31:0] r7541_out;
	wire [31:0] r7542_out;
	wire [31:0] r7543_out;
	wire [31:0] r7544_out;
	wire [31:0] r7545_out;
	wire [31:0] r7546_out;
	wire [31:0] r7547_out;
	wire [31:0] r7548_out;
	wire [31:0] r7549_out;
	wire [31:0] r7550_out;
	wire [31:0] r7551_out;
	wire [31:0] r7552_out;
	wire [31:0] r7553_out;
	wire [31:0] r7554_out;
	wire [31:0] r7555_out;
	wire [31:0] r7556_out;
	wire [31:0] r7557_out;
	wire [31:0] r7558_out;
	wire [31:0] r7559_out;
	wire [31:0] r7560_out;
	wire [31:0] r7561_out;
	wire [31:0] r7562_out;
	wire [31:0] r7563_out;
	wire [31:0] r7564_out;
	wire [31:0] r7565_out;
	wire [31:0] r7566_out;
	wire [31:0] r7567_out;
	wire [31:0] r7568_out;
	wire [31:0] r7569_out;
	wire [31:0] r7570_out;
	wire [31:0] r7571_out;
	wire [31:0] r7572_out;
	wire [31:0] r7573_out;
	wire [31:0] r7574_out;
	wire [31:0] r7575_out;
	wire [31:0] r7576_out;
	wire [31:0] r7577_out;
	wire [31:0] r7578_out;
	wire [31:0] r7579_out;
	wire [31:0] r7580_out;
	wire [31:0] r7581_out;
	wire [31:0] r7582_out;
	wire [31:0] r7583_out;
	wire [31:0] r7584_out;
	wire [31:0] r7585_out;
	wire [31:0] r7586_out;
	wire [31:0] r7587_out;
	wire [31:0] r7588_out;
	wire [31:0] r7589_out;
	wire [31:0] r7590_out;
	wire [31:0] r7591_out;
	wire [31:0] r7592_out;
	wire [31:0] r7593_out;
	wire [31:0] r7594_out;
	wire [31:0] r7595_out;
	wire [31:0] r7596_out;
	wire [31:0] r7597_out;
	wire [31:0] r7598_out;
	wire [31:0] r7599_out;
	wire [31:0] r7600_out;
	wire [31:0] r7601_out;
	wire [31:0] r7602_out;
	wire [31:0] r7603_out;
	wire [31:0] r7604_out;
	wire [31:0] r7605_out;
	wire [31:0] r7606_out;
	wire [31:0] r7607_out;
	wire [31:0] r7608_out;
	wire [31:0] r7609_out;
	wire [31:0] r7610_out;
	wire [31:0] r7611_out;
	wire [31:0] r7612_out;
	wire [31:0] r7613_out;
	wire [31:0] r7614_out;
	wire [31:0] r7615_out;
	wire [31:0] r7616_out;
	wire [31:0] r7617_out;
	wire [31:0] r7618_out;
	wire [31:0] r7619_out;
	wire [31:0] r7620_out;
	wire [31:0] r7621_out;
	wire [31:0] r7622_out;
	wire [31:0] r7623_out;
	wire [31:0] r7624_out;
	wire [31:0] r7625_out;
	wire [31:0] r7626_out;
	wire [31:0] r7627_out;
	wire [31:0] r7628_out;
	wire [31:0] r7629_out;
	wire [31:0] r7630_out;
	wire [31:0] r7631_out;
	wire [31:0] r7632_out;
	wire [31:0] r7633_out;
	wire [31:0] r7634_out;
	wire [31:0] r7635_out;
	wire [31:0] r7636_out;
	wire [31:0] r7637_out;
	wire [31:0] r7638_out;
	wire [31:0] r7639_out;
	wire [31:0] r7640_out;
	wire [31:0] r7641_out;
	wire [31:0] r7642_out;
	wire [31:0] r7643_out;
	wire [31:0] r7644_out;
	wire [31:0] r7645_out;
	wire [31:0] r7646_out;
	wire [31:0] r7647_out;
	wire [31:0] r7648_out;
	wire [31:0] r7649_out;
	wire [31:0] r7650_out;
	wire [31:0] r7651_out;
	wire [31:0] r7652_out;
	wire [31:0] r7653_out;
	wire [31:0] r7654_out;
	wire [31:0] r7655_out;
	wire [31:0] r7656_out;
	wire [31:0] r7657_out;
	wire [31:0] r7658_out;
	wire [31:0] r7659_out;
	wire [31:0] r7660_out;
	wire [31:0] r7661_out;
	wire [31:0] r7662_out;
	wire [31:0] r7663_out;
	wire [31:0] r7664_out;
	wire [31:0] r7665_out;
	wire [31:0] r7666_out;
	wire [31:0] r7667_out;
	wire [31:0] r7668_out;
	wire [31:0] r7669_out;
	wire [31:0] r7670_out;
	wire [31:0] r7671_out;
	wire [31:0] r7672_out;
	wire [31:0] r7673_out;
	wire [31:0] r7674_out;
	wire [31:0] r7675_out;
	wire [31:0] r7676_out;
	wire [31:0] r7677_out;
	wire [31:0] r7678_out;
	wire [31:0] r7679_out;
	wire [31:0] r7680_out;
	wire [31:0] r7681_out;
	wire [31:0] r7682_out;
	wire [31:0] r7683_out;
	wire [31:0] r7684_out;
	wire [31:0] r7685_out;
	wire [31:0] r7686_out;
	wire [31:0] r7687_out;
	wire [31:0] r7688_out;
	wire [31:0] r7689_out;
	wire [31:0] r7690_out;
	wire [31:0] r7691_out;
	wire [31:0] r7692_out;
	wire [31:0] r7693_out;
	wire [31:0] r7694_out;
	wire [31:0] r7695_out;
	wire [31:0] r7696_out;
	wire [31:0] r7697_out;
	wire [31:0] r7698_out;
	wire [31:0] r7699_out;
	wire [31:0] r7700_out;
	wire [31:0] r7701_out;
	wire [31:0] r7702_out;
	wire [31:0] r7703_out;
	wire [31:0] r7704_out;
	wire [31:0] r7705_out;
	wire [31:0] r7706_out;
	wire [31:0] r7707_out;
	wire [31:0] r7708_out;
	wire [31:0] r7709_out;
	wire [31:0] r7710_out;
	wire [31:0] r7711_out;
	wire [31:0] r7712_out;
	wire [31:0] r7713_out;
	wire [31:0] r7714_out;
	wire [31:0] r7715_out;
	wire [31:0] r7716_out;
	wire [31:0] r7717_out;
	wire [31:0] r7718_out;
	wire [31:0] r7719_out;
	wire [31:0] r7720_out;
	wire [31:0] r7721_out;
	wire [31:0] r7722_out;
	wire [31:0] r7723_out;
	wire [31:0] r7724_out;
	wire [31:0] r7725_out;
	wire [31:0] r7726_out;
	wire [31:0] r7727_out;
	wire [31:0] r7728_out;
	wire [31:0] r7729_out;
	wire [31:0] r7730_out;
	wire [31:0] r7731_out;
	wire [31:0] r7732_out;
	wire [31:0] r7733_out;
	wire [31:0] r7734_out;
	wire [31:0] r7735_out;
	wire [31:0] r7736_out;
	wire [31:0] r7737_out;
	wire [31:0] r7738_out;
	wire [31:0] r7739_out;
	wire [31:0] r7740_out;
	wire [31:0] r7741_out;
	wire [31:0] r7742_out;
	wire [31:0] r7743_out;
	wire [31:0] r7744_out;
	wire [31:0] r7745_out;
	wire [31:0] r7746_out;
	wire [31:0] r7747_out;
	wire [31:0] r7748_out;
	wire [31:0] r7749_out;
	wire [31:0] r7750_out;
	wire [31:0] r7751_out;
	wire [31:0] r7752_out;
	wire [31:0] r7753_out;
	wire [31:0] r7754_out;
	wire [31:0] r7755_out;
	wire [31:0] r7756_out;
	wire [31:0] r7757_out;
	wire [31:0] r7758_out;
	wire [31:0] r7759_out;
	wire [31:0] r7760_out;
	wire [31:0] r7761_out;
	wire [31:0] r7762_out;
	wire [31:0] r7763_out;
	wire [31:0] r7764_out;
	wire [31:0] r7765_out;
	wire [31:0] r7766_out;
	wire [31:0] r7767_out;
	wire [31:0] r7768_out;
	wire [31:0] r7769_out;
	wire [31:0] r7770_out;
	wire [31:0] r7771_out;
	wire [31:0] r7772_out;
	wire [31:0] r7773_out;
	wire [31:0] r7774_out;
	wire [31:0] r7775_out;
	wire [31:0] r7776_out;
	wire [31:0] r7777_out;
	wire [31:0] r7778_out;
	wire [31:0] r7779_out;
	wire [31:0] r7780_out;
	wire [31:0] r7781_out;
	wire [31:0] r7782_out;
	wire [31:0] r7783_out;
	wire [31:0] r7784_out;
	wire [31:0] r7785_out;
	wire [31:0] r7786_out;
	wire [31:0] r7787_out;
	wire [31:0] r7788_out;
	wire [31:0] r7789_out;
	wire [31:0] r7790_out;
	wire [31:0] r7791_out;
	wire [31:0] r7792_out;
	wire [31:0] r7793_out;
	wire [31:0] r7794_out;
	wire [31:0] r7795_out;
	wire [31:0] r7796_out;
	wire [31:0] r7797_out;
	wire [31:0] r7798_out;
	wire [31:0] r7799_out;
	wire [31:0] r7800_out;
	wire [31:0] r7801_out;
	wire [31:0] r7802_out;
	wire [31:0] r7803_out;
	wire [31:0] r7804_out;
	wire [31:0] r7805_out;
	wire [31:0] r7806_out;
	wire [31:0] r7807_out;
	wire [31:0] r7808_out;
	wire [31:0] r7809_out;
	wire [31:0] r7810_out;
	wire [31:0] r7811_out;
	wire [31:0] r7812_out;
	wire [31:0] r7813_out;
	wire [31:0] r7814_out;
	wire [31:0] r7815_out;
	wire [31:0] r7816_out;
	wire [31:0] r7817_out;
	wire [31:0] r7818_out;
	wire [31:0] r7819_out;
	wire [31:0] r7820_out;
	wire [31:0] r7821_out;
	wire [31:0] r7822_out;
	wire [31:0] r7823_out;
	wire [31:0] r7824_out;
	wire [31:0] r7825_out;
	wire [31:0] r7826_out;
	wire [31:0] r7827_out;
	wire [31:0] r7828_out;
	wire [31:0] r7829_out;
	wire [31:0] r7830_out;
	wire [31:0] r7831_out;
	wire [31:0] r7832_out;
	wire [31:0] r7833_out;
	wire [31:0] r7834_out;
	wire [31:0] r7835_out;
	wire [31:0] r7836_out;
	wire [31:0] r7837_out;
	wire [31:0] r7838_out;
	wire [31:0] r7839_out;
	wire [31:0] r7840_out;
	wire [31:0] r7841_out;
	wire [31:0] r7842_out;
	wire [31:0] r7843_out;
	wire [31:0] r7844_out;
	wire [31:0] r7845_out;
	wire [31:0] r7846_out;
	wire [31:0] r7847_out;
	wire [31:0] r7848_out;
	wire [31:0] r7849_out;
	wire [31:0] r7850_out;
	wire [31:0] r7851_out;
	wire [31:0] r7852_out;
	wire [31:0] r7853_out;
	wire [31:0] r7854_out;
	wire [31:0] r7855_out;
	wire [31:0] r7856_out;
	wire [31:0] r7857_out;
	wire [31:0] r7858_out;
	wire [31:0] r7859_out;
	wire [31:0] r7860_out;
	wire [31:0] r7861_out;
	wire [31:0] r7862_out;
	wire [31:0] r7863_out;
	wire [31:0] r7864_out;
	wire [31:0] r7865_out;
	wire [31:0] r7866_out;
	wire [31:0] r7867_out;
	wire [31:0] r7868_out;
	wire [31:0] r7869_out;
	wire [31:0] r7870_out;
	wire [31:0] r7871_out;
	wire [31:0] r7872_out;
	wire [31:0] r7873_out;
	wire [31:0] r7874_out;
	wire [31:0] r7875_out;
	wire [31:0] r7876_out;
	wire [31:0] r7877_out;
	wire [31:0] r7878_out;
	wire [31:0] r7879_out;
	wire [31:0] r7880_out;
	wire [31:0] r7881_out;
	wire [31:0] r7882_out;
	wire [31:0] r7883_out;
	wire [31:0] r7884_out;
	wire [31:0] r7885_out;
	wire [31:0] r7886_out;
	wire [31:0] r7887_out;
	wire [31:0] r7888_out;
	wire [31:0] r7889_out;
	wire [31:0] r7890_out;
	wire [31:0] r7891_out;
	wire [31:0] r7892_out;
	wire [31:0] r7893_out;
	wire [31:0] r7894_out;
	wire [31:0] r7895_out;
	wire [31:0] r7896_out;
	wire [31:0] r7897_out;
	wire [31:0] r7898_out;
	wire [31:0] r7899_out;
	wire [31:0] r7900_out;
	wire [31:0] r7901_out;
	wire [31:0] r7902_out;
	wire [31:0] r7903_out;
	wire [31:0] r7904_out;
	wire [31:0] r7905_out;
	wire [31:0] r7906_out;
	wire [31:0] r7907_out;
	wire [31:0] r7908_out;
	wire [31:0] r7909_out;
	wire [31:0] r7910_out;
	wire [31:0] r7911_out;
	wire [31:0] r7912_out;
	wire [31:0] r7913_out;
	wire [31:0] r7914_out;
	wire [31:0] r7915_out;
	wire [31:0] r7916_out;
	wire [31:0] r7917_out;
	wire [31:0] r7918_out;
	wire [31:0] r7919_out;
	wire [31:0] r7920_out;
	wire [31:0] r7921_out;
	wire [31:0] r7922_out;
	wire [31:0] r7923_out;
	wire [31:0] r7924_out;
	wire [31:0] r7925_out;
	wire [31:0] r7926_out;
	wire [31:0] r7927_out;
	wire [31:0] r7928_out;
	wire [31:0] r7929_out;
	wire [31:0] r7930_out;
	wire [31:0] r7931_out;
	wire [31:0] r7932_out;
	wire [31:0] r7933_out;
	wire [31:0] r7934_out;
	wire [31:0] r7935_out;
	wire [31:0] r7936_out;
	wire [31:0] r7937_out;
	wire [31:0] r7938_out;
	wire [31:0] r7939_out;
	wire [31:0] r7940_out;
	wire [31:0] r7941_out;
	wire [31:0] r7942_out;
	wire [31:0] r7943_out;
	wire [31:0] r7944_out;
	wire [31:0] r7945_out;
	wire [31:0] r7946_out;
	wire [31:0] r7947_out;
	wire [31:0] r7948_out;
	wire [31:0] r7949_out;
	wire [31:0] r7950_out;
	wire [31:0] r7951_out;
	wire [31:0] r7952_out;
	wire [31:0] r7953_out;
	wire [31:0] r7954_out;
	wire [31:0] r7955_out;
	wire [31:0] r7956_out;
	wire [31:0] r7957_out;
	wire [31:0] r7958_out;
	wire [31:0] r7959_out;
	wire [31:0] r7960_out;
	wire [31:0] r7961_out;
	wire [31:0] r7962_out;
	wire [31:0] r7963_out;
	wire [31:0] r7964_out;
	wire [31:0] r7965_out;
	wire [31:0] r7966_out;
	wire [31:0] r7967_out;
	wire [31:0] r7968_out;
	wire [31:0] r7969_out;
	wire [31:0] r7970_out;
	wire [31:0] r7971_out;
	wire [31:0] r7972_out;
	wire [31:0] r7973_out;
	wire [31:0] r7974_out;
	wire [31:0] r7975_out;
	wire [31:0] r7976_out;
	wire [31:0] r7977_out;
	wire [31:0] r7978_out;
	wire [31:0] r7979_out;
	wire [31:0] r7980_out;
	wire [31:0] r7981_out;
	wire [31:0] r7982_out;
	wire [31:0] r7983_out;
	wire [31:0] r7984_out;
	wire [31:0] r7985_out;
	wire [31:0] r7986_out;
	wire [31:0] r7987_out;
	wire [31:0] r7988_out;
	wire [31:0] r7989_out;
	wire [31:0] r7990_out;
	wire [31:0] r7991_out;
	wire [31:0] r7992_out;
	wire [31:0] r7993_out;
	wire [31:0] r7994_out;
	wire [31:0] r7995_out;
	wire [31:0] r7996_out;
	wire [31:0] r7997_out;
	wire [31:0] r7998_out;
	wire [31:0] r7999_out;

	reg32 r0 (rst, clk, in, r0_out);
	reg32 r1 (rst, clk, in, r1_out);
	reg32 r2 (rst, clk, in, r2_out);
	reg32 r3 (rst, clk, in, r3_out);
	reg32 r4 (rst, clk, in, r4_out);
	reg32 r5 (rst, clk, in, r5_out);
	reg32 r6 (rst, clk, in, r6_out);
	reg32 r7 (rst, clk, in, r7_out);
	reg32 r8 (rst, clk, in, r8_out);
	reg32 r9 (rst, clk, in, r9_out);
	reg32 r10 (rst, clk, in, r10_out);
	reg32 r11 (rst, clk, in, r11_out);
	reg32 r12 (rst, clk, in, r12_out);
	reg32 r13 (rst, clk, in, r13_out);
	reg32 r14 (rst, clk, in, r14_out);
	reg32 r15 (rst, clk, in, r15_out);
	reg32 r16 (rst, clk, in, r16_out);
	reg32 r17 (rst, clk, in, r17_out);
	reg32 r18 (rst, clk, in, r18_out);
	reg32 r19 (rst, clk, in, r19_out);
	reg32 r20 (rst, clk, in, r20_out);
	reg32 r21 (rst, clk, in, r21_out);
	reg32 r22 (rst, clk, in, r22_out);
	reg32 r23 (rst, clk, in, r23_out);
	reg32 r24 (rst, clk, in, r24_out);
	reg32 r25 (rst, clk, in, r25_out);
	reg32 r26 (rst, clk, in, r26_out);
	reg32 r27 (rst, clk, in, r27_out);
	reg32 r28 (rst, clk, in, r28_out);
	reg32 r29 (rst, clk, in, r29_out);
	reg32 r30 (rst, clk, in, r30_out);
	reg32 r31 (rst, clk, in, r31_out);
	reg32 r32 (rst, clk, in, r32_out);
	reg32 r33 (rst, clk, in, r33_out);
	reg32 r34 (rst, clk, in, r34_out);
	reg32 r35 (rst, clk, in, r35_out);
	reg32 r36 (rst, clk, in, r36_out);
	reg32 r37 (rst, clk, in, r37_out);
	reg32 r38 (rst, clk, in, r38_out);
	reg32 r39 (rst, clk, in, r39_out);
	reg32 r40 (rst, clk, in, r40_out);
	reg32 r41 (rst, clk, in, r41_out);
	reg32 r42 (rst, clk, in, r42_out);
	reg32 r43 (rst, clk, in, r43_out);
	reg32 r44 (rst, clk, in, r44_out);
	reg32 r45 (rst, clk, in, r45_out);
	reg32 r46 (rst, clk, in, r46_out);
	reg32 r47 (rst, clk, in, r47_out);
	reg32 r48 (rst, clk, in, r48_out);
	reg32 r49 (rst, clk, in, r49_out);
	reg32 r50 (rst, clk, in, r50_out);
	reg32 r51 (rst, clk, in, r51_out);
	reg32 r52 (rst, clk, in, r52_out);
	reg32 r53 (rst, clk, in, r53_out);
	reg32 r54 (rst, clk, in, r54_out);
	reg32 r55 (rst, clk, in, r55_out);
	reg32 r56 (rst, clk, in, r56_out);
	reg32 r57 (rst, clk, in, r57_out);
	reg32 r58 (rst, clk, in, r58_out);
	reg32 r59 (rst, clk, in, r59_out);
	reg32 r60 (rst, clk, in, r60_out);
	reg32 r61 (rst, clk, in, r61_out);
	reg32 r62 (rst, clk, in, r62_out);
	reg32 r63 (rst, clk, in, r63_out);
	reg32 r64 (rst, clk, in, r64_out);
	reg32 r65 (rst, clk, in, r65_out);
	reg32 r66 (rst, clk, in, r66_out);
	reg32 r67 (rst, clk, in, r67_out);
	reg32 r68 (rst, clk, in, r68_out);
	reg32 r69 (rst, clk, in, r69_out);
	reg32 r70 (rst, clk, in, r70_out);
	reg32 r71 (rst, clk, in, r71_out);
	reg32 r72 (rst, clk, in, r72_out);
	reg32 r73 (rst, clk, in, r73_out);
	reg32 r74 (rst, clk, in, r74_out);
	reg32 r75 (rst, clk, in, r75_out);
	reg32 r76 (rst, clk, in, r76_out);
	reg32 r77 (rst, clk, in, r77_out);
	reg32 r78 (rst, clk, in, r78_out);
	reg32 r79 (rst, clk, in, r79_out);
	reg32 r80 (rst, clk, in, r80_out);
	reg32 r81 (rst, clk, in, r81_out);
	reg32 r82 (rst, clk, in, r82_out);
	reg32 r83 (rst, clk, in, r83_out);
	reg32 r84 (rst, clk, in, r84_out);
	reg32 r85 (rst, clk, in, r85_out);
	reg32 r86 (rst, clk, in, r86_out);
	reg32 r87 (rst, clk, in, r87_out);
	reg32 r88 (rst, clk, in, r88_out);
	reg32 r89 (rst, clk, in, r89_out);
	reg32 r90 (rst, clk, in, r90_out);
	reg32 r91 (rst, clk, in, r91_out);
	reg32 r92 (rst, clk, in, r92_out);
	reg32 r93 (rst, clk, in, r93_out);
	reg32 r94 (rst, clk, in, r94_out);
	reg32 r95 (rst, clk, in, r95_out);
	reg32 r96 (rst, clk, in, r96_out);
	reg32 r97 (rst, clk, in, r97_out);
	reg32 r98 (rst, clk, in, r98_out);
	reg32 r99 (rst, clk, in, r99_out);
	reg32 r100 (rst, clk, in, r100_out);
	reg32 r101 (rst, clk, in, r101_out);
	reg32 r102 (rst, clk, in, r102_out);
	reg32 r103 (rst, clk, in, r103_out);
	reg32 r104 (rst, clk, in, r104_out);
	reg32 r105 (rst, clk, in, r105_out);
	reg32 r106 (rst, clk, in, r106_out);
	reg32 r107 (rst, clk, in, r107_out);
	reg32 r108 (rst, clk, in, r108_out);
	reg32 r109 (rst, clk, in, r109_out);
	reg32 r110 (rst, clk, in, r110_out);
	reg32 r111 (rst, clk, in, r111_out);
	reg32 r112 (rst, clk, in, r112_out);
	reg32 r113 (rst, clk, in, r113_out);
	reg32 r114 (rst, clk, in, r114_out);
	reg32 r115 (rst, clk, in, r115_out);
	reg32 r116 (rst, clk, in, r116_out);
	reg32 r117 (rst, clk, in, r117_out);
	reg32 r118 (rst, clk, in, r118_out);
	reg32 r119 (rst, clk, in, r119_out);
	reg32 r120 (rst, clk, in, r120_out);
	reg32 r121 (rst, clk, in, r121_out);
	reg32 r122 (rst, clk, in, r122_out);
	reg32 r123 (rst, clk, in, r123_out);
	reg32 r124 (rst, clk, in, r124_out);
	reg32 r125 (rst, clk, in, r125_out);
	reg32 r126 (rst, clk, in, r126_out);
	reg32 r127 (rst, clk, in, r127_out);
	reg32 r128 (rst, clk, in, r128_out);
	reg32 r129 (rst, clk, in, r129_out);
	reg32 r130 (rst, clk, in, r130_out);
	reg32 r131 (rst, clk, in, r131_out);
	reg32 r132 (rst, clk, in, r132_out);
	reg32 r133 (rst, clk, in, r133_out);
	reg32 r134 (rst, clk, in, r134_out);
	reg32 r135 (rst, clk, in, r135_out);
	reg32 r136 (rst, clk, in, r136_out);
	reg32 r137 (rst, clk, in, r137_out);
	reg32 r138 (rst, clk, in, r138_out);
	reg32 r139 (rst, clk, in, r139_out);
	reg32 r140 (rst, clk, in, r140_out);
	reg32 r141 (rst, clk, in, r141_out);
	reg32 r142 (rst, clk, in, r142_out);
	reg32 r143 (rst, clk, in, r143_out);
	reg32 r144 (rst, clk, in, r144_out);
	reg32 r145 (rst, clk, in, r145_out);
	reg32 r146 (rst, clk, in, r146_out);
	reg32 r147 (rst, clk, in, r147_out);
	reg32 r148 (rst, clk, in, r148_out);
	reg32 r149 (rst, clk, in, r149_out);
	reg32 r150 (rst, clk, in, r150_out);
	reg32 r151 (rst, clk, in, r151_out);
	reg32 r152 (rst, clk, in, r152_out);
	reg32 r153 (rst, clk, in, r153_out);
	reg32 r154 (rst, clk, in, r154_out);
	reg32 r155 (rst, clk, in, r155_out);
	reg32 r156 (rst, clk, in, r156_out);
	reg32 r157 (rst, clk, in, r157_out);
	reg32 r158 (rst, clk, in, r158_out);
	reg32 r159 (rst, clk, in, r159_out);
	reg32 r160 (rst, clk, in, r160_out);
	reg32 r161 (rst, clk, in, r161_out);
	reg32 r162 (rst, clk, in, r162_out);
	reg32 r163 (rst, clk, in, r163_out);
	reg32 r164 (rst, clk, in, r164_out);
	reg32 r165 (rst, clk, in, r165_out);
	reg32 r166 (rst, clk, in, r166_out);
	reg32 r167 (rst, clk, in, r167_out);
	reg32 r168 (rst, clk, in, r168_out);
	reg32 r169 (rst, clk, in, r169_out);
	reg32 r170 (rst, clk, in, r170_out);
	reg32 r171 (rst, clk, in, r171_out);
	reg32 r172 (rst, clk, in, r172_out);
	reg32 r173 (rst, clk, in, r173_out);
	reg32 r174 (rst, clk, in, r174_out);
	reg32 r175 (rst, clk, in, r175_out);
	reg32 r176 (rst, clk, in, r176_out);
	reg32 r177 (rst, clk, in, r177_out);
	reg32 r178 (rst, clk, in, r178_out);
	reg32 r179 (rst, clk, in, r179_out);
	reg32 r180 (rst, clk, in, r180_out);
	reg32 r181 (rst, clk, in, r181_out);
	reg32 r182 (rst, clk, in, r182_out);
	reg32 r183 (rst, clk, in, r183_out);
	reg32 r184 (rst, clk, in, r184_out);
	reg32 r185 (rst, clk, in, r185_out);
	reg32 r186 (rst, clk, in, r186_out);
	reg32 r187 (rst, clk, in, r187_out);
	reg32 r188 (rst, clk, in, r188_out);
	reg32 r189 (rst, clk, in, r189_out);
	reg32 r190 (rst, clk, in, r190_out);
	reg32 r191 (rst, clk, in, r191_out);
	reg32 r192 (rst, clk, in, r192_out);
	reg32 r193 (rst, clk, in, r193_out);
	reg32 r194 (rst, clk, in, r194_out);
	reg32 r195 (rst, clk, in, r195_out);
	reg32 r196 (rst, clk, in, r196_out);
	reg32 r197 (rst, clk, in, r197_out);
	reg32 r198 (rst, clk, in, r198_out);
	reg32 r199 (rst, clk, in, r199_out);
	reg32 r200 (rst, clk, in, r200_out);
	reg32 r201 (rst, clk, in, r201_out);
	reg32 r202 (rst, clk, in, r202_out);
	reg32 r203 (rst, clk, in, r203_out);
	reg32 r204 (rst, clk, in, r204_out);
	reg32 r205 (rst, clk, in, r205_out);
	reg32 r206 (rst, clk, in, r206_out);
	reg32 r207 (rst, clk, in, r207_out);
	reg32 r208 (rst, clk, in, r208_out);
	reg32 r209 (rst, clk, in, r209_out);
	reg32 r210 (rst, clk, in, r210_out);
	reg32 r211 (rst, clk, in, r211_out);
	reg32 r212 (rst, clk, in, r212_out);
	reg32 r213 (rst, clk, in, r213_out);
	reg32 r214 (rst, clk, in, r214_out);
	reg32 r215 (rst, clk, in, r215_out);
	reg32 r216 (rst, clk, in, r216_out);
	reg32 r217 (rst, clk, in, r217_out);
	reg32 r218 (rst, clk, in, r218_out);
	reg32 r219 (rst, clk, in, r219_out);
	reg32 r220 (rst, clk, in, r220_out);
	reg32 r221 (rst, clk, in, r221_out);
	reg32 r222 (rst, clk, in, r222_out);
	reg32 r223 (rst, clk, in, r223_out);
	reg32 r224 (rst, clk, in, r224_out);
	reg32 r225 (rst, clk, in, r225_out);
	reg32 r226 (rst, clk, in, r226_out);
	reg32 r227 (rst, clk, in, r227_out);
	reg32 r228 (rst, clk, in, r228_out);
	reg32 r229 (rst, clk, in, r229_out);
	reg32 r230 (rst, clk, in, r230_out);
	reg32 r231 (rst, clk, in, r231_out);
	reg32 r232 (rst, clk, in, r232_out);
	reg32 r233 (rst, clk, in, r233_out);
	reg32 r234 (rst, clk, in, r234_out);
	reg32 r235 (rst, clk, in, r235_out);
	reg32 r236 (rst, clk, in, r236_out);
	reg32 r237 (rst, clk, in, r237_out);
	reg32 r238 (rst, clk, in, r238_out);
	reg32 r239 (rst, clk, in, r239_out);
	reg32 r240 (rst, clk, in, r240_out);
	reg32 r241 (rst, clk, in, r241_out);
	reg32 r242 (rst, clk, in, r242_out);
	reg32 r243 (rst, clk, in, r243_out);
	reg32 r244 (rst, clk, in, r244_out);
	reg32 r245 (rst, clk, in, r245_out);
	reg32 r246 (rst, clk, in, r246_out);
	reg32 r247 (rst, clk, in, r247_out);
	reg32 r248 (rst, clk, in, r248_out);
	reg32 r249 (rst, clk, in, r249_out);
	reg32 r250 (rst, clk, in, r250_out);
	reg32 r251 (rst, clk, in, r251_out);
	reg32 r252 (rst, clk, in, r252_out);
	reg32 r253 (rst, clk, in, r253_out);
	reg32 r254 (rst, clk, in, r254_out);
	reg32 r255 (rst, clk, in, r255_out);
	reg32 r256 (rst, clk, in, r256_out);
	reg32 r257 (rst, clk, in, r257_out);
	reg32 r258 (rst, clk, in, r258_out);
	reg32 r259 (rst, clk, in, r259_out);
	reg32 r260 (rst, clk, in, r260_out);
	reg32 r261 (rst, clk, in, r261_out);
	reg32 r262 (rst, clk, in, r262_out);
	reg32 r263 (rst, clk, in, r263_out);
	reg32 r264 (rst, clk, in, r264_out);
	reg32 r265 (rst, clk, in, r265_out);
	reg32 r266 (rst, clk, in, r266_out);
	reg32 r267 (rst, clk, in, r267_out);
	reg32 r268 (rst, clk, in, r268_out);
	reg32 r269 (rst, clk, in, r269_out);
	reg32 r270 (rst, clk, in, r270_out);
	reg32 r271 (rst, clk, in, r271_out);
	reg32 r272 (rst, clk, in, r272_out);
	reg32 r273 (rst, clk, in, r273_out);
	reg32 r274 (rst, clk, in, r274_out);
	reg32 r275 (rst, clk, in, r275_out);
	reg32 r276 (rst, clk, in, r276_out);
	reg32 r277 (rst, clk, in, r277_out);
	reg32 r278 (rst, clk, in, r278_out);
	reg32 r279 (rst, clk, in, r279_out);
	reg32 r280 (rst, clk, in, r280_out);
	reg32 r281 (rst, clk, in, r281_out);
	reg32 r282 (rst, clk, in, r282_out);
	reg32 r283 (rst, clk, in, r283_out);
	reg32 r284 (rst, clk, in, r284_out);
	reg32 r285 (rst, clk, in, r285_out);
	reg32 r286 (rst, clk, in, r286_out);
	reg32 r287 (rst, clk, in, r287_out);
	reg32 r288 (rst, clk, in, r288_out);
	reg32 r289 (rst, clk, in, r289_out);
	reg32 r290 (rst, clk, in, r290_out);
	reg32 r291 (rst, clk, in, r291_out);
	reg32 r292 (rst, clk, in, r292_out);
	reg32 r293 (rst, clk, in, r293_out);
	reg32 r294 (rst, clk, in, r294_out);
	reg32 r295 (rst, clk, in, r295_out);
	reg32 r296 (rst, clk, in, r296_out);
	reg32 r297 (rst, clk, in, r297_out);
	reg32 r298 (rst, clk, in, r298_out);
	reg32 r299 (rst, clk, in, r299_out);
	reg32 r300 (rst, clk, in, r300_out);
	reg32 r301 (rst, clk, in, r301_out);
	reg32 r302 (rst, clk, in, r302_out);
	reg32 r303 (rst, clk, in, r303_out);
	reg32 r304 (rst, clk, in, r304_out);
	reg32 r305 (rst, clk, in, r305_out);
	reg32 r306 (rst, clk, in, r306_out);
	reg32 r307 (rst, clk, in, r307_out);
	reg32 r308 (rst, clk, in, r308_out);
	reg32 r309 (rst, clk, in, r309_out);
	reg32 r310 (rst, clk, in, r310_out);
	reg32 r311 (rst, clk, in, r311_out);
	reg32 r312 (rst, clk, in, r312_out);
	reg32 r313 (rst, clk, in, r313_out);
	reg32 r314 (rst, clk, in, r314_out);
	reg32 r315 (rst, clk, in, r315_out);
	reg32 r316 (rst, clk, in, r316_out);
	reg32 r317 (rst, clk, in, r317_out);
	reg32 r318 (rst, clk, in, r318_out);
	reg32 r319 (rst, clk, in, r319_out);
	reg32 r320 (rst, clk, in, r320_out);
	reg32 r321 (rst, clk, in, r321_out);
	reg32 r322 (rst, clk, in, r322_out);
	reg32 r323 (rst, clk, in, r323_out);
	reg32 r324 (rst, clk, in, r324_out);
	reg32 r325 (rst, clk, in, r325_out);
	reg32 r326 (rst, clk, in, r326_out);
	reg32 r327 (rst, clk, in, r327_out);
	reg32 r328 (rst, clk, in, r328_out);
	reg32 r329 (rst, clk, in, r329_out);
	reg32 r330 (rst, clk, in, r330_out);
	reg32 r331 (rst, clk, in, r331_out);
	reg32 r332 (rst, clk, in, r332_out);
	reg32 r333 (rst, clk, in, r333_out);
	reg32 r334 (rst, clk, in, r334_out);
	reg32 r335 (rst, clk, in, r335_out);
	reg32 r336 (rst, clk, in, r336_out);
	reg32 r337 (rst, clk, in, r337_out);
	reg32 r338 (rst, clk, in, r338_out);
	reg32 r339 (rst, clk, in, r339_out);
	reg32 r340 (rst, clk, in, r340_out);
	reg32 r341 (rst, clk, in, r341_out);
	reg32 r342 (rst, clk, in, r342_out);
	reg32 r343 (rst, clk, in, r343_out);
	reg32 r344 (rst, clk, in, r344_out);
	reg32 r345 (rst, clk, in, r345_out);
	reg32 r346 (rst, clk, in, r346_out);
	reg32 r347 (rst, clk, in, r347_out);
	reg32 r348 (rst, clk, in, r348_out);
	reg32 r349 (rst, clk, in, r349_out);
	reg32 r350 (rst, clk, in, r350_out);
	reg32 r351 (rst, clk, in, r351_out);
	reg32 r352 (rst, clk, in, r352_out);
	reg32 r353 (rst, clk, in, r353_out);
	reg32 r354 (rst, clk, in, r354_out);
	reg32 r355 (rst, clk, in, r355_out);
	reg32 r356 (rst, clk, in, r356_out);
	reg32 r357 (rst, clk, in, r357_out);
	reg32 r358 (rst, clk, in, r358_out);
	reg32 r359 (rst, clk, in, r359_out);
	reg32 r360 (rst, clk, in, r360_out);
	reg32 r361 (rst, clk, in, r361_out);
	reg32 r362 (rst, clk, in, r362_out);
	reg32 r363 (rst, clk, in, r363_out);
	reg32 r364 (rst, clk, in, r364_out);
	reg32 r365 (rst, clk, in, r365_out);
	reg32 r366 (rst, clk, in, r366_out);
	reg32 r367 (rst, clk, in, r367_out);
	reg32 r368 (rst, clk, in, r368_out);
	reg32 r369 (rst, clk, in, r369_out);
	reg32 r370 (rst, clk, in, r370_out);
	reg32 r371 (rst, clk, in, r371_out);
	reg32 r372 (rst, clk, in, r372_out);
	reg32 r373 (rst, clk, in, r373_out);
	reg32 r374 (rst, clk, in, r374_out);
	reg32 r375 (rst, clk, in, r375_out);
	reg32 r376 (rst, clk, in, r376_out);
	reg32 r377 (rst, clk, in, r377_out);
	reg32 r378 (rst, clk, in, r378_out);
	reg32 r379 (rst, clk, in, r379_out);
	reg32 r380 (rst, clk, in, r380_out);
	reg32 r381 (rst, clk, in, r381_out);
	reg32 r382 (rst, clk, in, r382_out);
	reg32 r383 (rst, clk, in, r383_out);
	reg32 r384 (rst, clk, in, r384_out);
	reg32 r385 (rst, clk, in, r385_out);
	reg32 r386 (rst, clk, in, r386_out);
	reg32 r387 (rst, clk, in, r387_out);
	reg32 r388 (rst, clk, in, r388_out);
	reg32 r389 (rst, clk, in, r389_out);
	reg32 r390 (rst, clk, in, r390_out);
	reg32 r391 (rst, clk, in, r391_out);
	reg32 r392 (rst, clk, in, r392_out);
	reg32 r393 (rst, clk, in, r393_out);
	reg32 r394 (rst, clk, in, r394_out);
	reg32 r395 (rst, clk, in, r395_out);
	reg32 r396 (rst, clk, in, r396_out);
	reg32 r397 (rst, clk, in, r397_out);
	reg32 r398 (rst, clk, in, r398_out);
	reg32 r399 (rst, clk, in, r399_out);
	reg32 r400 (rst, clk, in, r400_out);
	reg32 r401 (rst, clk, in, r401_out);
	reg32 r402 (rst, clk, in, r402_out);
	reg32 r403 (rst, clk, in, r403_out);
	reg32 r404 (rst, clk, in, r404_out);
	reg32 r405 (rst, clk, in, r405_out);
	reg32 r406 (rst, clk, in, r406_out);
	reg32 r407 (rst, clk, in, r407_out);
	reg32 r408 (rst, clk, in, r408_out);
	reg32 r409 (rst, clk, in, r409_out);
	reg32 r410 (rst, clk, in, r410_out);
	reg32 r411 (rst, clk, in, r411_out);
	reg32 r412 (rst, clk, in, r412_out);
	reg32 r413 (rst, clk, in, r413_out);
	reg32 r414 (rst, clk, in, r414_out);
	reg32 r415 (rst, clk, in, r415_out);
	reg32 r416 (rst, clk, in, r416_out);
	reg32 r417 (rst, clk, in, r417_out);
	reg32 r418 (rst, clk, in, r418_out);
	reg32 r419 (rst, clk, in, r419_out);
	reg32 r420 (rst, clk, in, r420_out);
	reg32 r421 (rst, clk, in, r421_out);
	reg32 r422 (rst, clk, in, r422_out);
	reg32 r423 (rst, clk, in, r423_out);
	reg32 r424 (rst, clk, in, r424_out);
	reg32 r425 (rst, clk, in, r425_out);
	reg32 r426 (rst, clk, in, r426_out);
	reg32 r427 (rst, clk, in, r427_out);
	reg32 r428 (rst, clk, in, r428_out);
	reg32 r429 (rst, clk, in, r429_out);
	reg32 r430 (rst, clk, in, r430_out);
	reg32 r431 (rst, clk, in, r431_out);
	reg32 r432 (rst, clk, in, r432_out);
	reg32 r433 (rst, clk, in, r433_out);
	reg32 r434 (rst, clk, in, r434_out);
	reg32 r435 (rst, clk, in, r435_out);
	reg32 r436 (rst, clk, in, r436_out);
	reg32 r437 (rst, clk, in, r437_out);
	reg32 r438 (rst, clk, in, r438_out);
	reg32 r439 (rst, clk, in, r439_out);
	reg32 r440 (rst, clk, in, r440_out);
	reg32 r441 (rst, clk, in, r441_out);
	reg32 r442 (rst, clk, in, r442_out);
	reg32 r443 (rst, clk, in, r443_out);
	reg32 r444 (rst, clk, in, r444_out);
	reg32 r445 (rst, clk, in, r445_out);
	reg32 r446 (rst, clk, in, r446_out);
	reg32 r447 (rst, clk, in, r447_out);
	reg32 r448 (rst, clk, in, r448_out);
	reg32 r449 (rst, clk, in, r449_out);
	reg32 r450 (rst, clk, in, r450_out);
	reg32 r451 (rst, clk, in, r451_out);
	reg32 r452 (rst, clk, in, r452_out);
	reg32 r453 (rst, clk, in, r453_out);
	reg32 r454 (rst, clk, in, r454_out);
	reg32 r455 (rst, clk, in, r455_out);
	reg32 r456 (rst, clk, in, r456_out);
	reg32 r457 (rst, clk, in, r457_out);
	reg32 r458 (rst, clk, in, r458_out);
	reg32 r459 (rst, clk, in, r459_out);
	reg32 r460 (rst, clk, in, r460_out);
	reg32 r461 (rst, clk, in, r461_out);
	reg32 r462 (rst, clk, in, r462_out);
	reg32 r463 (rst, clk, in, r463_out);
	reg32 r464 (rst, clk, in, r464_out);
	reg32 r465 (rst, clk, in, r465_out);
	reg32 r466 (rst, clk, in, r466_out);
	reg32 r467 (rst, clk, in, r467_out);
	reg32 r468 (rst, clk, in, r468_out);
	reg32 r469 (rst, clk, in, r469_out);
	reg32 r470 (rst, clk, in, r470_out);
	reg32 r471 (rst, clk, in, r471_out);
	reg32 r472 (rst, clk, in, r472_out);
	reg32 r473 (rst, clk, in, r473_out);
	reg32 r474 (rst, clk, in, r474_out);
	reg32 r475 (rst, clk, in, r475_out);
	reg32 r476 (rst, clk, in, r476_out);
	reg32 r477 (rst, clk, in, r477_out);
	reg32 r478 (rst, clk, in, r478_out);
	reg32 r479 (rst, clk, in, r479_out);
	reg32 r480 (rst, clk, in, r480_out);
	reg32 r481 (rst, clk, in, r481_out);
	reg32 r482 (rst, clk, in, r482_out);
	reg32 r483 (rst, clk, in, r483_out);
	reg32 r484 (rst, clk, in, r484_out);
	reg32 r485 (rst, clk, in, r485_out);
	reg32 r486 (rst, clk, in, r486_out);
	reg32 r487 (rst, clk, in, r487_out);
	reg32 r488 (rst, clk, in, r488_out);
	reg32 r489 (rst, clk, in, r489_out);
	reg32 r490 (rst, clk, in, r490_out);
	reg32 r491 (rst, clk, in, r491_out);
	reg32 r492 (rst, clk, in, r492_out);
	reg32 r493 (rst, clk, in, r493_out);
	reg32 r494 (rst, clk, in, r494_out);
	reg32 r495 (rst, clk, in, r495_out);
	reg32 r496 (rst, clk, in, r496_out);
	reg32 r497 (rst, clk, in, r497_out);
	reg32 r498 (rst, clk, in, r498_out);
	reg32 r499 (rst, clk, in, r499_out);
	reg32 r500 (rst, clk, in, r500_out);
	reg32 r501 (rst, clk, in, r501_out);
	reg32 r502 (rst, clk, in, r502_out);
	reg32 r503 (rst, clk, in, r503_out);
	reg32 r504 (rst, clk, in, r504_out);
	reg32 r505 (rst, clk, in, r505_out);
	reg32 r506 (rst, clk, in, r506_out);
	reg32 r507 (rst, clk, in, r507_out);
	reg32 r508 (rst, clk, in, r508_out);
	reg32 r509 (rst, clk, in, r509_out);
	reg32 r510 (rst, clk, in, r510_out);
	reg32 r511 (rst, clk, in, r511_out);
	reg32 r512 (rst, clk, in, r512_out);
	reg32 r513 (rst, clk, in, r513_out);
	reg32 r514 (rst, clk, in, r514_out);
	reg32 r515 (rst, clk, in, r515_out);
	reg32 r516 (rst, clk, in, r516_out);
	reg32 r517 (rst, clk, in, r517_out);
	reg32 r518 (rst, clk, in, r518_out);
	reg32 r519 (rst, clk, in, r519_out);
	reg32 r520 (rst, clk, in, r520_out);
	reg32 r521 (rst, clk, in, r521_out);
	reg32 r522 (rst, clk, in, r522_out);
	reg32 r523 (rst, clk, in, r523_out);
	reg32 r524 (rst, clk, in, r524_out);
	reg32 r525 (rst, clk, in, r525_out);
	reg32 r526 (rst, clk, in, r526_out);
	reg32 r527 (rst, clk, in, r527_out);
	reg32 r528 (rst, clk, in, r528_out);
	reg32 r529 (rst, clk, in, r529_out);
	reg32 r530 (rst, clk, in, r530_out);
	reg32 r531 (rst, clk, in, r531_out);
	reg32 r532 (rst, clk, in, r532_out);
	reg32 r533 (rst, clk, in, r533_out);
	reg32 r534 (rst, clk, in, r534_out);
	reg32 r535 (rst, clk, in, r535_out);
	reg32 r536 (rst, clk, in, r536_out);
	reg32 r537 (rst, clk, in, r537_out);
	reg32 r538 (rst, clk, in, r538_out);
	reg32 r539 (rst, clk, in, r539_out);
	reg32 r540 (rst, clk, in, r540_out);
	reg32 r541 (rst, clk, in, r541_out);
	reg32 r542 (rst, clk, in, r542_out);
	reg32 r543 (rst, clk, in, r543_out);
	reg32 r544 (rst, clk, in, r544_out);
	reg32 r545 (rst, clk, in, r545_out);
	reg32 r546 (rst, clk, in, r546_out);
	reg32 r547 (rst, clk, in, r547_out);
	reg32 r548 (rst, clk, in, r548_out);
	reg32 r549 (rst, clk, in, r549_out);
	reg32 r550 (rst, clk, in, r550_out);
	reg32 r551 (rst, clk, in, r551_out);
	reg32 r552 (rst, clk, in, r552_out);
	reg32 r553 (rst, clk, in, r553_out);
	reg32 r554 (rst, clk, in, r554_out);
	reg32 r555 (rst, clk, in, r555_out);
	reg32 r556 (rst, clk, in, r556_out);
	reg32 r557 (rst, clk, in, r557_out);
	reg32 r558 (rst, clk, in, r558_out);
	reg32 r559 (rst, clk, in, r559_out);
	reg32 r560 (rst, clk, in, r560_out);
	reg32 r561 (rst, clk, in, r561_out);
	reg32 r562 (rst, clk, in, r562_out);
	reg32 r563 (rst, clk, in, r563_out);
	reg32 r564 (rst, clk, in, r564_out);
	reg32 r565 (rst, clk, in, r565_out);
	reg32 r566 (rst, clk, in, r566_out);
	reg32 r567 (rst, clk, in, r567_out);
	reg32 r568 (rst, clk, in, r568_out);
	reg32 r569 (rst, clk, in, r569_out);
	reg32 r570 (rst, clk, in, r570_out);
	reg32 r571 (rst, clk, in, r571_out);
	reg32 r572 (rst, clk, in, r572_out);
	reg32 r573 (rst, clk, in, r573_out);
	reg32 r574 (rst, clk, in, r574_out);
	reg32 r575 (rst, clk, in, r575_out);
	reg32 r576 (rst, clk, in, r576_out);
	reg32 r577 (rst, clk, in, r577_out);
	reg32 r578 (rst, clk, in, r578_out);
	reg32 r579 (rst, clk, in, r579_out);
	reg32 r580 (rst, clk, in, r580_out);
	reg32 r581 (rst, clk, in, r581_out);
	reg32 r582 (rst, clk, in, r582_out);
	reg32 r583 (rst, clk, in, r583_out);
	reg32 r584 (rst, clk, in, r584_out);
	reg32 r585 (rst, clk, in, r585_out);
	reg32 r586 (rst, clk, in, r586_out);
	reg32 r587 (rst, clk, in, r587_out);
	reg32 r588 (rst, clk, in, r588_out);
	reg32 r589 (rst, clk, in, r589_out);
	reg32 r590 (rst, clk, in, r590_out);
	reg32 r591 (rst, clk, in, r591_out);
	reg32 r592 (rst, clk, in, r592_out);
	reg32 r593 (rst, clk, in, r593_out);
	reg32 r594 (rst, clk, in, r594_out);
	reg32 r595 (rst, clk, in, r595_out);
	reg32 r596 (rst, clk, in, r596_out);
	reg32 r597 (rst, clk, in, r597_out);
	reg32 r598 (rst, clk, in, r598_out);
	reg32 r599 (rst, clk, in, r599_out);
	reg32 r600 (rst, clk, in, r600_out);
	reg32 r601 (rst, clk, in, r601_out);
	reg32 r602 (rst, clk, in, r602_out);
	reg32 r603 (rst, clk, in, r603_out);
	reg32 r604 (rst, clk, in, r604_out);
	reg32 r605 (rst, clk, in, r605_out);
	reg32 r606 (rst, clk, in, r606_out);
	reg32 r607 (rst, clk, in, r607_out);
	reg32 r608 (rst, clk, in, r608_out);
	reg32 r609 (rst, clk, in, r609_out);
	reg32 r610 (rst, clk, in, r610_out);
	reg32 r611 (rst, clk, in, r611_out);
	reg32 r612 (rst, clk, in, r612_out);
	reg32 r613 (rst, clk, in, r613_out);
	reg32 r614 (rst, clk, in, r614_out);
	reg32 r615 (rst, clk, in, r615_out);
	reg32 r616 (rst, clk, in, r616_out);
	reg32 r617 (rst, clk, in, r617_out);
	reg32 r618 (rst, clk, in, r618_out);
	reg32 r619 (rst, clk, in, r619_out);
	reg32 r620 (rst, clk, in, r620_out);
	reg32 r621 (rst, clk, in, r621_out);
	reg32 r622 (rst, clk, in, r622_out);
	reg32 r623 (rst, clk, in, r623_out);
	reg32 r624 (rst, clk, in, r624_out);
	reg32 r625 (rst, clk, in, r625_out);
	reg32 r626 (rst, clk, in, r626_out);
	reg32 r627 (rst, clk, in, r627_out);
	reg32 r628 (rst, clk, in, r628_out);
	reg32 r629 (rst, clk, in, r629_out);
	reg32 r630 (rst, clk, in, r630_out);
	reg32 r631 (rst, clk, in, r631_out);
	reg32 r632 (rst, clk, in, r632_out);
	reg32 r633 (rst, clk, in, r633_out);
	reg32 r634 (rst, clk, in, r634_out);
	reg32 r635 (rst, clk, in, r635_out);
	reg32 r636 (rst, clk, in, r636_out);
	reg32 r637 (rst, clk, in, r637_out);
	reg32 r638 (rst, clk, in, r638_out);
	reg32 r639 (rst, clk, in, r639_out);
	reg32 r640 (rst, clk, in, r640_out);
	reg32 r641 (rst, clk, in, r641_out);
	reg32 r642 (rst, clk, in, r642_out);
	reg32 r643 (rst, clk, in, r643_out);
	reg32 r644 (rst, clk, in, r644_out);
	reg32 r645 (rst, clk, in, r645_out);
	reg32 r646 (rst, clk, in, r646_out);
	reg32 r647 (rst, clk, in, r647_out);
	reg32 r648 (rst, clk, in, r648_out);
	reg32 r649 (rst, clk, in, r649_out);
	reg32 r650 (rst, clk, in, r650_out);
	reg32 r651 (rst, clk, in, r651_out);
	reg32 r652 (rst, clk, in, r652_out);
	reg32 r653 (rst, clk, in, r653_out);
	reg32 r654 (rst, clk, in, r654_out);
	reg32 r655 (rst, clk, in, r655_out);
	reg32 r656 (rst, clk, in, r656_out);
	reg32 r657 (rst, clk, in, r657_out);
	reg32 r658 (rst, clk, in, r658_out);
	reg32 r659 (rst, clk, in, r659_out);
	reg32 r660 (rst, clk, in, r660_out);
	reg32 r661 (rst, clk, in, r661_out);
	reg32 r662 (rst, clk, in, r662_out);
	reg32 r663 (rst, clk, in, r663_out);
	reg32 r664 (rst, clk, in, r664_out);
	reg32 r665 (rst, clk, in, r665_out);
	reg32 r666 (rst, clk, in, r666_out);
	reg32 r667 (rst, clk, in, r667_out);
	reg32 r668 (rst, clk, in, r668_out);
	reg32 r669 (rst, clk, in, r669_out);
	reg32 r670 (rst, clk, in, r670_out);
	reg32 r671 (rst, clk, in, r671_out);
	reg32 r672 (rst, clk, in, r672_out);
	reg32 r673 (rst, clk, in, r673_out);
	reg32 r674 (rst, clk, in, r674_out);
	reg32 r675 (rst, clk, in, r675_out);
	reg32 r676 (rst, clk, in, r676_out);
	reg32 r677 (rst, clk, in, r677_out);
	reg32 r678 (rst, clk, in, r678_out);
	reg32 r679 (rst, clk, in, r679_out);
	reg32 r680 (rst, clk, in, r680_out);
	reg32 r681 (rst, clk, in, r681_out);
	reg32 r682 (rst, clk, in, r682_out);
	reg32 r683 (rst, clk, in, r683_out);
	reg32 r684 (rst, clk, in, r684_out);
	reg32 r685 (rst, clk, in, r685_out);
	reg32 r686 (rst, clk, in, r686_out);
	reg32 r687 (rst, clk, in, r687_out);
	reg32 r688 (rst, clk, in, r688_out);
	reg32 r689 (rst, clk, in, r689_out);
	reg32 r690 (rst, clk, in, r690_out);
	reg32 r691 (rst, clk, in, r691_out);
	reg32 r692 (rst, clk, in, r692_out);
	reg32 r693 (rst, clk, in, r693_out);
	reg32 r694 (rst, clk, in, r694_out);
	reg32 r695 (rst, clk, in, r695_out);
	reg32 r696 (rst, clk, in, r696_out);
	reg32 r697 (rst, clk, in, r697_out);
	reg32 r698 (rst, clk, in, r698_out);
	reg32 r699 (rst, clk, in, r699_out);
	reg32 r700 (rst, clk, in, r700_out);
	reg32 r701 (rst, clk, in, r701_out);
	reg32 r702 (rst, clk, in, r702_out);
	reg32 r703 (rst, clk, in, r703_out);
	reg32 r704 (rst, clk, in, r704_out);
	reg32 r705 (rst, clk, in, r705_out);
	reg32 r706 (rst, clk, in, r706_out);
	reg32 r707 (rst, clk, in, r707_out);
	reg32 r708 (rst, clk, in, r708_out);
	reg32 r709 (rst, clk, in, r709_out);
	reg32 r710 (rst, clk, in, r710_out);
	reg32 r711 (rst, clk, in, r711_out);
	reg32 r712 (rst, clk, in, r712_out);
	reg32 r713 (rst, clk, in, r713_out);
	reg32 r714 (rst, clk, in, r714_out);
	reg32 r715 (rst, clk, in, r715_out);
	reg32 r716 (rst, clk, in, r716_out);
	reg32 r717 (rst, clk, in, r717_out);
	reg32 r718 (rst, clk, in, r718_out);
	reg32 r719 (rst, clk, in, r719_out);
	reg32 r720 (rst, clk, in, r720_out);
	reg32 r721 (rst, clk, in, r721_out);
	reg32 r722 (rst, clk, in, r722_out);
	reg32 r723 (rst, clk, in, r723_out);
	reg32 r724 (rst, clk, in, r724_out);
	reg32 r725 (rst, clk, in, r725_out);
	reg32 r726 (rst, clk, in, r726_out);
	reg32 r727 (rst, clk, in, r727_out);
	reg32 r728 (rst, clk, in, r728_out);
	reg32 r729 (rst, clk, in, r729_out);
	reg32 r730 (rst, clk, in, r730_out);
	reg32 r731 (rst, clk, in, r731_out);
	reg32 r732 (rst, clk, in, r732_out);
	reg32 r733 (rst, clk, in, r733_out);
	reg32 r734 (rst, clk, in, r734_out);
	reg32 r735 (rst, clk, in, r735_out);
	reg32 r736 (rst, clk, in, r736_out);
	reg32 r737 (rst, clk, in, r737_out);
	reg32 r738 (rst, clk, in, r738_out);
	reg32 r739 (rst, clk, in, r739_out);
	reg32 r740 (rst, clk, in, r740_out);
	reg32 r741 (rst, clk, in, r741_out);
	reg32 r742 (rst, clk, in, r742_out);
	reg32 r743 (rst, clk, in, r743_out);
	reg32 r744 (rst, clk, in, r744_out);
	reg32 r745 (rst, clk, in, r745_out);
	reg32 r746 (rst, clk, in, r746_out);
	reg32 r747 (rst, clk, in, r747_out);
	reg32 r748 (rst, clk, in, r748_out);
	reg32 r749 (rst, clk, in, r749_out);
	reg32 r750 (rst, clk, in, r750_out);
	reg32 r751 (rst, clk, in, r751_out);
	reg32 r752 (rst, clk, in, r752_out);
	reg32 r753 (rst, clk, in, r753_out);
	reg32 r754 (rst, clk, in, r754_out);
	reg32 r755 (rst, clk, in, r755_out);
	reg32 r756 (rst, clk, in, r756_out);
	reg32 r757 (rst, clk, in, r757_out);
	reg32 r758 (rst, clk, in, r758_out);
	reg32 r759 (rst, clk, in, r759_out);
	reg32 r760 (rst, clk, in, r760_out);
	reg32 r761 (rst, clk, in, r761_out);
	reg32 r762 (rst, clk, in, r762_out);
	reg32 r763 (rst, clk, in, r763_out);
	reg32 r764 (rst, clk, in, r764_out);
	reg32 r765 (rst, clk, in, r765_out);
	reg32 r766 (rst, clk, in, r766_out);
	reg32 r767 (rst, clk, in, r767_out);
	reg32 r768 (rst, clk, in, r768_out);
	reg32 r769 (rst, clk, in, r769_out);
	reg32 r770 (rst, clk, in, r770_out);
	reg32 r771 (rst, clk, in, r771_out);
	reg32 r772 (rst, clk, in, r772_out);
	reg32 r773 (rst, clk, in, r773_out);
	reg32 r774 (rst, clk, in, r774_out);
	reg32 r775 (rst, clk, in, r775_out);
	reg32 r776 (rst, clk, in, r776_out);
	reg32 r777 (rst, clk, in, r777_out);
	reg32 r778 (rst, clk, in, r778_out);
	reg32 r779 (rst, clk, in, r779_out);
	reg32 r780 (rst, clk, in, r780_out);
	reg32 r781 (rst, clk, in, r781_out);
	reg32 r782 (rst, clk, in, r782_out);
	reg32 r783 (rst, clk, in, r783_out);
	reg32 r784 (rst, clk, in, r784_out);
	reg32 r785 (rst, clk, in, r785_out);
	reg32 r786 (rst, clk, in, r786_out);
	reg32 r787 (rst, clk, in, r787_out);
	reg32 r788 (rst, clk, in, r788_out);
	reg32 r789 (rst, clk, in, r789_out);
	reg32 r790 (rst, clk, in, r790_out);
	reg32 r791 (rst, clk, in, r791_out);
	reg32 r792 (rst, clk, in, r792_out);
	reg32 r793 (rst, clk, in, r793_out);
	reg32 r794 (rst, clk, in, r794_out);
	reg32 r795 (rst, clk, in, r795_out);
	reg32 r796 (rst, clk, in, r796_out);
	reg32 r797 (rst, clk, in, r797_out);
	reg32 r798 (rst, clk, in, r798_out);
	reg32 r799 (rst, clk, in, r799_out);
	reg32 r800 (rst, clk, in, r800_out);
	reg32 r801 (rst, clk, in, r801_out);
	reg32 r802 (rst, clk, in, r802_out);
	reg32 r803 (rst, clk, in, r803_out);
	reg32 r804 (rst, clk, in, r804_out);
	reg32 r805 (rst, clk, in, r805_out);
	reg32 r806 (rst, clk, in, r806_out);
	reg32 r807 (rst, clk, in, r807_out);
	reg32 r808 (rst, clk, in, r808_out);
	reg32 r809 (rst, clk, in, r809_out);
	reg32 r810 (rst, clk, in, r810_out);
	reg32 r811 (rst, clk, in, r811_out);
	reg32 r812 (rst, clk, in, r812_out);
	reg32 r813 (rst, clk, in, r813_out);
	reg32 r814 (rst, clk, in, r814_out);
	reg32 r815 (rst, clk, in, r815_out);
	reg32 r816 (rst, clk, in, r816_out);
	reg32 r817 (rst, clk, in, r817_out);
	reg32 r818 (rst, clk, in, r818_out);
	reg32 r819 (rst, clk, in, r819_out);
	reg32 r820 (rst, clk, in, r820_out);
	reg32 r821 (rst, clk, in, r821_out);
	reg32 r822 (rst, clk, in, r822_out);
	reg32 r823 (rst, clk, in, r823_out);
	reg32 r824 (rst, clk, in, r824_out);
	reg32 r825 (rst, clk, in, r825_out);
	reg32 r826 (rst, clk, in, r826_out);
	reg32 r827 (rst, clk, in, r827_out);
	reg32 r828 (rst, clk, in, r828_out);
	reg32 r829 (rst, clk, in, r829_out);
	reg32 r830 (rst, clk, in, r830_out);
	reg32 r831 (rst, clk, in, r831_out);
	reg32 r832 (rst, clk, in, r832_out);
	reg32 r833 (rst, clk, in, r833_out);
	reg32 r834 (rst, clk, in, r834_out);
	reg32 r835 (rst, clk, in, r835_out);
	reg32 r836 (rst, clk, in, r836_out);
	reg32 r837 (rst, clk, in, r837_out);
	reg32 r838 (rst, clk, in, r838_out);
	reg32 r839 (rst, clk, in, r839_out);
	reg32 r840 (rst, clk, in, r840_out);
	reg32 r841 (rst, clk, in, r841_out);
	reg32 r842 (rst, clk, in, r842_out);
	reg32 r843 (rst, clk, in, r843_out);
	reg32 r844 (rst, clk, in, r844_out);
	reg32 r845 (rst, clk, in, r845_out);
	reg32 r846 (rst, clk, in, r846_out);
	reg32 r847 (rst, clk, in, r847_out);
	reg32 r848 (rst, clk, in, r848_out);
	reg32 r849 (rst, clk, in, r849_out);
	reg32 r850 (rst, clk, in, r850_out);
	reg32 r851 (rst, clk, in, r851_out);
	reg32 r852 (rst, clk, in, r852_out);
	reg32 r853 (rst, clk, in, r853_out);
	reg32 r854 (rst, clk, in, r854_out);
	reg32 r855 (rst, clk, in, r855_out);
	reg32 r856 (rst, clk, in, r856_out);
	reg32 r857 (rst, clk, in, r857_out);
	reg32 r858 (rst, clk, in, r858_out);
	reg32 r859 (rst, clk, in, r859_out);
	reg32 r860 (rst, clk, in, r860_out);
	reg32 r861 (rst, clk, in, r861_out);
	reg32 r862 (rst, clk, in, r862_out);
	reg32 r863 (rst, clk, in, r863_out);
	reg32 r864 (rst, clk, in, r864_out);
	reg32 r865 (rst, clk, in, r865_out);
	reg32 r866 (rst, clk, in, r866_out);
	reg32 r867 (rst, clk, in, r867_out);
	reg32 r868 (rst, clk, in, r868_out);
	reg32 r869 (rst, clk, in, r869_out);
	reg32 r870 (rst, clk, in, r870_out);
	reg32 r871 (rst, clk, in, r871_out);
	reg32 r872 (rst, clk, in, r872_out);
	reg32 r873 (rst, clk, in, r873_out);
	reg32 r874 (rst, clk, in, r874_out);
	reg32 r875 (rst, clk, in, r875_out);
	reg32 r876 (rst, clk, in, r876_out);
	reg32 r877 (rst, clk, in, r877_out);
	reg32 r878 (rst, clk, in, r878_out);
	reg32 r879 (rst, clk, in, r879_out);
	reg32 r880 (rst, clk, in, r880_out);
	reg32 r881 (rst, clk, in, r881_out);
	reg32 r882 (rst, clk, in, r882_out);
	reg32 r883 (rst, clk, in, r883_out);
	reg32 r884 (rst, clk, in, r884_out);
	reg32 r885 (rst, clk, in, r885_out);
	reg32 r886 (rst, clk, in, r886_out);
	reg32 r887 (rst, clk, in, r887_out);
	reg32 r888 (rst, clk, in, r888_out);
	reg32 r889 (rst, clk, in, r889_out);
	reg32 r890 (rst, clk, in, r890_out);
	reg32 r891 (rst, clk, in, r891_out);
	reg32 r892 (rst, clk, in, r892_out);
	reg32 r893 (rst, clk, in, r893_out);
	reg32 r894 (rst, clk, in, r894_out);
	reg32 r895 (rst, clk, in, r895_out);
	reg32 r896 (rst, clk, in, r896_out);
	reg32 r897 (rst, clk, in, r897_out);
	reg32 r898 (rst, clk, in, r898_out);
	reg32 r899 (rst, clk, in, r899_out);
	reg32 r900 (rst, clk, in, r900_out);
	reg32 r901 (rst, clk, in, r901_out);
	reg32 r902 (rst, clk, in, r902_out);
	reg32 r903 (rst, clk, in, r903_out);
	reg32 r904 (rst, clk, in, r904_out);
	reg32 r905 (rst, clk, in, r905_out);
	reg32 r906 (rst, clk, in, r906_out);
	reg32 r907 (rst, clk, in, r907_out);
	reg32 r908 (rst, clk, in, r908_out);
	reg32 r909 (rst, clk, in, r909_out);
	reg32 r910 (rst, clk, in, r910_out);
	reg32 r911 (rst, clk, in, r911_out);
	reg32 r912 (rst, clk, in, r912_out);
	reg32 r913 (rst, clk, in, r913_out);
	reg32 r914 (rst, clk, in, r914_out);
	reg32 r915 (rst, clk, in, r915_out);
	reg32 r916 (rst, clk, in, r916_out);
	reg32 r917 (rst, clk, in, r917_out);
	reg32 r918 (rst, clk, in, r918_out);
	reg32 r919 (rst, clk, in, r919_out);
	reg32 r920 (rst, clk, in, r920_out);
	reg32 r921 (rst, clk, in, r921_out);
	reg32 r922 (rst, clk, in, r922_out);
	reg32 r923 (rst, clk, in, r923_out);
	reg32 r924 (rst, clk, in, r924_out);
	reg32 r925 (rst, clk, in, r925_out);
	reg32 r926 (rst, clk, in, r926_out);
	reg32 r927 (rst, clk, in, r927_out);
	reg32 r928 (rst, clk, in, r928_out);
	reg32 r929 (rst, clk, in, r929_out);
	reg32 r930 (rst, clk, in, r930_out);
	reg32 r931 (rst, clk, in, r931_out);
	reg32 r932 (rst, clk, in, r932_out);
	reg32 r933 (rst, clk, in, r933_out);
	reg32 r934 (rst, clk, in, r934_out);
	reg32 r935 (rst, clk, in, r935_out);
	reg32 r936 (rst, clk, in, r936_out);
	reg32 r937 (rst, clk, in, r937_out);
	reg32 r938 (rst, clk, in, r938_out);
	reg32 r939 (rst, clk, in, r939_out);
	reg32 r940 (rst, clk, in, r940_out);
	reg32 r941 (rst, clk, in, r941_out);
	reg32 r942 (rst, clk, in, r942_out);
	reg32 r943 (rst, clk, in, r943_out);
	reg32 r944 (rst, clk, in, r944_out);
	reg32 r945 (rst, clk, in, r945_out);
	reg32 r946 (rst, clk, in, r946_out);
	reg32 r947 (rst, clk, in, r947_out);
	reg32 r948 (rst, clk, in, r948_out);
	reg32 r949 (rst, clk, in, r949_out);
	reg32 r950 (rst, clk, in, r950_out);
	reg32 r951 (rst, clk, in, r951_out);
	reg32 r952 (rst, clk, in, r952_out);
	reg32 r953 (rst, clk, in, r953_out);
	reg32 r954 (rst, clk, in, r954_out);
	reg32 r955 (rst, clk, in, r955_out);
	reg32 r956 (rst, clk, in, r956_out);
	reg32 r957 (rst, clk, in, r957_out);
	reg32 r958 (rst, clk, in, r958_out);
	reg32 r959 (rst, clk, in, r959_out);
	reg32 r960 (rst, clk, in, r960_out);
	reg32 r961 (rst, clk, in, r961_out);
	reg32 r962 (rst, clk, in, r962_out);
	reg32 r963 (rst, clk, in, r963_out);
	reg32 r964 (rst, clk, in, r964_out);
	reg32 r965 (rst, clk, in, r965_out);
	reg32 r966 (rst, clk, in, r966_out);
	reg32 r967 (rst, clk, in, r967_out);
	reg32 r968 (rst, clk, in, r968_out);
	reg32 r969 (rst, clk, in, r969_out);
	reg32 r970 (rst, clk, in, r970_out);
	reg32 r971 (rst, clk, in, r971_out);
	reg32 r972 (rst, clk, in, r972_out);
	reg32 r973 (rst, clk, in, r973_out);
	reg32 r974 (rst, clk, in, r974_out);
	reg32 r975 (rst, clk, in, r975_out);
	reg32 r976 (rst, clk, in, r976_out);
	reg32 r977 (rst, clk, in, r977_out);
	reg32 r978 (rst, clk, in, r978_out);
	reg32 r979 (rst, clk, in, r979_out);
	reg32 r980 (rst, clk, in, r980_out);
	reg32 r981 (rst, clk, in, r981_out);
	reg32 r982 (rst, clk, in, r982_out);
	reg32 r983 (rst, clk, in, r983_out);
	reg32 r984 (rst, clk, in, r984_out);
	reg32 r985 (rst, clk, in, r985_out);
	reg32 r986 (rst, clk, in, r986_out);
	reg32 r987 (rst, clk, in, r987_out);
	reg32 r988 (rst, clk, in, r988_out);
	reg32 r989 (rst, clk, in, r989_out);
	reg32 r990 (rst, clk, in, r990_out);
	reg32 r991 (rst, clk, in, r991_out);
	reg32 r992 (rst, clk, in, r992_out);
	reg32 r993 (rst, clk, in, r993_out);
	reg32 r994 (rst, clk, in, r994_out);
	reg32 r995 (rst, clk, in, r995_out);
	reg32 r996 (rst, clk, in, r996_out);
	reg32 r997 (rst, clk, in, r997_out);
	reg32 r998 (rst, clk, in, r998_out);
	reg32 r999 (rst, clk, in, r999_out);
	reg32 r1000 (rst, clk, in, r1000_out);
	reg32 r1001 (rst, clk, in, r1001_out);
	reg32 r1002 (rst, clk, in, r1002_out);
	reg32 r1003 (rst, clk, in, r1003_out);
	reg32 r1004 (rst, clk, in, r1004_out);
	reg32 r1005 (rst, clk, in, r1005_out);
	reg32 r1006 (rst, clk, in, r1006_out);
	reg32 r1007 (rst, clk, in, r1007_out);
	reg32 r1008 (rst, clk, in, r1008_out);
	reg32 r1009 (rst, clk, in, r1009_out);
	reg32 r1010 (rst, clk, in, r1010_out);
	reg32 r1011 (rst, clk, in, r1011_out);
	reg32 r1012 (rst, clk, in, r1012_out);
	reg32 r1013 (rst, clk, in, r1013_out);
	reg32 r1014 (rst, clk, in, r1014_out);
	reg32 r1015 (rst, clk, in, r1015_out);
	reg32 r1016 (rst, clk, in, r1016_out);
	reg32 r1017 (rst, clk, in, r1017_out);
	reg32 r1018 (rst, clk, in, r1018_out);
	reg32 r1019 (rst, clk, in, r1019_out);
	reg32 r1020 (rst, clk, in, r1020_out);
	reg32 r1021 (rst, clk, in, r1021_out);
	reg32 r1022 (rst, clk, in, r1022_out);
	reg32 r1023 (rst, clk, in, r1023_out);
	reg32 r1024 (rst, clk, in, r1024_out);
	reg32 r1025 (rst, clk, in, r1025_out);
	reg32 r1026 (rst, clk, in, r1026_out);
	reg32 r1027 (rst, clk, in, r1027_out);
	reg32 r1028 (rst, clk, in, r1028_out);
	reg32 r1029 (rst, clk, in, r1029_out);
	reg32 r1030 (rst, clk, in, r1030_out);
	reg32 r1031 (rst, clk, in, r1031_out);
	reg32 r1032 (rst, clk, in, r1032_out);
	reg32 r1033 (rst, clk, in, r1033_out);
	reg32 r1034 (rst, clk, in, r1034_out);
	reg32 r1035 (rst, clk, in, r1035_out);
	reg32 r1036 (rst, clk, in, r1036_out);
	reg32 r1037 (rst, clk, in, r1037_out);
	reg32 r1038 (rst, clk, in, r1038_out);
	reg32 r1039 (rst, clk, in, r1039_out);
	reg32 r1040 (rst, clk, in, r1040_out);
	reg32 r1041 (rst, clk, in, r1041_out);
	reg32 r1042 (rst, clk, in, r1042_out);
	reg32 r1043 (rst, clk, in, r1043_out);
	reg32 r1044 (rst, clk, in, r1044_out);
	reg32 r1045 (rst, clk, in, r1045_out);
	reg32 r1046 (rst, clk, in, r1046_out);
	reg32 r1047 (rst, clk, in, r1047_out);
	reg32 r1048 (rst, clk, in, r1048_out);
	reg32 r1049 (rst, clk, in, r1049_out);
	reg32 r1050 (rst, clk, in, r1050_out);
	reg32 r1051 (rst, clk, in, r1051_out);
	reg32 r1052 (rst, clk, in, r1052_out);
	reg32 r1053 (rst, clk, in, r1053_out);
	reg32 r1054 (rst, clk, in, r1054_out);
	reg32 r1055 (rst, clk, in, r1055_out);
	reg32 r1056 (rst, clk, in, r1056_out);
	reg32 r1057 (rst, clk, in, r1057_out);
	reg32 r1058 (rst, clk, in, r1058_out);
	reg32 r1059 (rst, clk, in, r1059_out);
	reg32 r1060 (rst, clk, in, r1060_out);
	reg32 r1061 (rst, clk, in, r1061_out);
	reg32 r1062 (rst, clk, in, r1062_out);
	reg32 r1063 (rst, clk, in, r1063_out);
	reg32 r1064 (rst, clk, in, r1064_out);
	reg32 r1065 (rst, clk, in, r1065_out);
	reg32 r1066 (rst, clk, in, r1066_out);
	reg32 r1067 (rst, clk, in, r1067_out);
	reg32 r1068 (rst, clk, in, r1068_out);
	reg32 r1069 (rst, clk, in, r1069_out);
	reg32 r1070 (rst, clk, in, r1070_out);
	reg32 r1071 (rst, clk, in, r1071_out);
	reg32 r1072 (rst, clk, in, r1072_out);
	reg32 r1073 (rst, clk, in, r1073_out);
	reg32 r1074 (rst, clk, in, r1074_out);
	reg32 r1075 (rst, clk, in, r1075_out);
	reg32 r1076 (rst, clk, in, r1076_out);
	reg32 r1077 (rst, clk, in, r1077_out);
	reg32 r1078 (rst, clk, in, r1078_out);
	reg32 r1079 (rst, clk, in, r1079_out);
	reg32 r1080 (rst, clk, in, r1080_out);
	reg32 r1081 (rst, clk, in, r1081_out);
	reg32 r1082 (rst, clk, in, r1082_out);
	reg32 r1083 (rst, clk, in, r1083_out);
	reg32 r1084 (rst, clk, in, r1084_out);
	reg32 r1085 (rst, clk, in, r1085_out);
	reg32 r1086 (rst, clk, in, r1086_out);
	reg32 r1087 (rst, clk, in, r1087_out);
	reg32 r1088 (rst, clk, in, r1088_out);
	reg32 r1089 (rst, clk, in, r1089_out);
	reg32 r1090 (rst, clk, in, r1090_out);
	reg32 r1091 (rst, clk, in, r1091_out);
	reg32 r1092 (rst, clk, in, r1092_out);
	reg32 r1093 (rst, clk, in, r1093_out);
	reg32 r1094 (rst, clk, in, r1094_out);
	reg32 r1095 (rst, clk, in, r1095_out);
	reg32 r1096 (rst, clk, in, r1096_out);
	reg32 r1097 (rst, clk, in, r1097_out);
	reg32 r1098 (rst, clk, in, r1098_out);
	reg32 r1099 (rst, clk, in, r1099_out);
	reg32 r1100 (rst, clk, in, r1100_out);
	reg32 r1101 (rst, clk, in, r1101_out);
	reg32 r1102 (rst, clk, in, r1102_out);
	reg32 r1103 (rst, clk, in, r1103_out);
	reg32 r1104 (rst, clk, in, r1104_out);
	reg32 r1105 (rst, clk, in, r1105_out);
	reg32 r1106 (rst, clk, in, r1106_out);
	reg32 r1107 (rst, clk, in, r1107_out);
	reg32 r1108 (rst, clk, in, r1108_out);
	reg32 r1109 (rst, clk, in, r1109_out);
	reg32 r1110 (rst, clk, in, r1110_out);
	reg32 r1111 (rst, clk, in, r1111_out);
	reg32 r1112 (rst, clk, in, r1112_out);
	reg32 r1113 (rst, clk, in, r1113_out);
	reg32 r1114 (rst, clk, in, r1114_out);
	reg32 r1115 (rst, clk, in, r1115_out);
	reg32 r1116 (rst, clk, in, r1116_out);
	reg32 r1117 (rst, clk, in, r1117_out);
	reg32 r1118 (rst, clk, in, r1118_out);
	reg32 r1119 (rst, clk, in, r1119_out);
	reg32 r1120 (rst, clk, in, r1120_out);
	reg32 r1121 (rst, clk, in, r1121_out);
	reg32 r1122 (rst, clk, in, r1122_out);
	reg32 r1123 (rst, clk, in, r1123_out);
	reg32 r1124 (rst, clk, in, r1124_out);
	reg32 r1125 (rst, clk, in, r1125_out);
	reg32 r1126 (rst, clk, in, r1126_out);
	reg32 r1127 (rst, clk, in, r1127_out);
	reg32 r1128 (rst, clk, in, r1128_out);
	reg32 r1129 (rst, clk, in, r1129_out);
	reg32 r1130 (rst, clk, in, r1130_out);
	reg32 r1131 (rst, clk, in, r1131_out);
	reg32 r1132 (rst, clk, in, r1132_out);
	reg32 r1133 (rst, clk, in, r1133_out);
	reg32 r1134 (rst, clk, in, r1134_out);
	reg32 r1135 (rst, clk, in, r1135_out);
	reg32 r1136 (rst, clk, in, r1136_out);
	reg32 r1137 (rst, clk, in, r1137_out);
	reg32 r1138 (rst, clk, in, r1138_out);
	reg32 r1139 (rst, clk, in, r1139_out);
	reg32 r1140 (rst, clk, in, r1140_out);
	reg32 r1141 (rst, clk, in, r1141_out);
	reg32 r1142 (rst, clk, in, r1142_out);
	reg32 r1143 (rst, clk, in, r1143_out);
	reg32 r1144 (rst, clk, in, r1144_out);
	reg32 r1145 (rst, clk, in, r1145_out);
	reg32 r1146 (rst, clk, in, r1146_out);
	reg32 r1147 (rst, clk, in, r1147_out);
	reg32 r1148 (rst, clk, in, r1148_out);
	reg32 r1149 (rst, clk, in, r1149_out);
	reg32 r1150 (rst, clk, in, r1150_out);
	reg32 r1151 (rst, clk, in, r1151_out);
	reg32 r1152 (rst, clk, in, r1152_out);
	reg32 r1153 (rst, clk, in, r1153_out);
	reg32 r1154 (rst, clk, in, r1154_out);
	reg32 r1155 (rst, clk, in, r1155_out);
	reg32 r1156 (rst, clk, in, r1156_out);
	reg32 r1157 (rst, clk, in, r1157_out);
	reg32 r1158 (rst, clk, in, r1158_out);
	reg32 r1159 (rst, clk, in, r1159_out);
	reg32 r1160 (rst, clk, in, r1160_out);
	reg32 r1161 (rst, clk, in, r1161_out);
	reg32 r1162 (rst, clk, in, r1162_out);
	reg32 r1163 (rst, clk, in, r1163_out);
	reg32 r1164 (rst, clk, in, r1164_out);
	reg32 r1165 (rst, clk, in, r1165_out);
	reg32 r1166 (rst, clk, in, r1166_out);
	reg32 r1167 (rst, clk, in, r1167_out);
	reg32 r1168 (rst, clk, in, r1168_out);
	reg32 r1169 (rst, clk, in, r1169_out);
	reg32 r1170 (rst, clk, in, r1170_out);
	reg32 r1171 (rst, clk, in, r1171_out);
	reg32 r1172 (rst, clk, in, r1172_out);
	reg32 r1173 (rst, clk, in, r1173_out);
	reg32 r1174 (rst, clk, in, r1174_out);
	reg32 r1175 (rst, clk, in, r1175_out);
	reg32 r1176 (rst, clk, in, r1176_out);
	reg32 r1177 (rst, clk, in, r1177_out);
	reg32 r1178 (rst, clk, in, r1178_out);
	reg32 r1179 (rst, clk, in, r1179_out);
	reg32 r1180 (rst, clk, in, r1180_out);
	reg32 r1181 (rst, clk, in, r1181_out);
	reg32 r1182 (rst, clk, in, r1182_out);
	reg32 r1183 (rst, clk, in, r1183_out);
	reg32 r1184 (rst, clk, in, r1184_out);
	reg32 r1185 (rst, clk, in, r1185_out);
	reg32 r1186 (rst, clk, in, r1186_out);
	reg32 r1187 (rst, clk, in, r1187_out);
	reg32 r1188 (rst, clk, in, r1188_out);
	reg32 r1189 (rst, clk, in, r1189_out);
	reg32 r1190 (rst, clk, in, r1190_out);
	reg32 r1191 (rst, clk, in, r1191_out);
	reg32 r1192 (rst, clk, in, r1192_out);
	reg32 r1193 (rst, clk, in, r1193_out);
	reg32 r1194 (rst, clk, in, r1194_out);
	reg32 r1195 (rst, clk, in, r1195_out);
	reg32 r1196 (rst, clk, in, r1196_out);
	reg32 r1197 (rst, clk, in, r1197_out);
	reg32 r1198 (rst, clk, in, r1198_out);
	reg32 r1199 (rst, clk, in, r1199_out);
	reg32 r1200 (rst, clk, in, r1200_out);
	reg32 r1201 (rst, clk, in, r1201_out);
	reg32 r1202 (rst, clk, in, r1202_out);
	reg32 r1203 (rst, clk, in, r1203_out);
	reg32 r1204 (rst, clk, in, r1204_out);
	reg32 r1205 (rst, clk, in, r1205_out);
	reg32 r1206 (rst, clk, in, r1206_out);
	reg32 r1207 (rst, clk, in, r1207_out);
	reg32 r1208 (rst, clk, in, r1208_out);
	reg32 r1209 (rst, clk, in, r1209_out);
	reg32 r1210 (rst, clk, in, r1210_out);
	reg32 r1211 (rst, clk, in, r1211_out);
	reg32 r1212 (rst, clk, in, r1212_out);
	reg32 r1213 (rst, clk, in, r1213_out);
	reg32 r1214 (rst, clk, in, r1214_out);
	reg32 r1215 (rst, clk, in, r1215_out);
	reg32 r1216 (rst, clk, in, r1216_out);
	reg32 r1217 (rst, clk, in, r1217_out);
	reg32 r1218 (rst, clk, in, r1218_out);
	reg32 r1219 (rst, clk, in, r1219_out);
	reg32 r1220 (rst, clk, in, r1220_out);
	reg32 r1221 (rst, clk, in, r1221_out);
	reg32 r1222 (rst, clk, in, r1222_out);
	reg32 r1223 (rst, clk, in, r1223_out);
	reg32 r1224 (rst, clk, in, r1224_out);
	reg32 r1225 (rst, clk, in, r1225_out);
	reg32 r1226 (rst, clk, in, r1226_out);
	reg32 r1227 (rst, clk, in, r1227_out);
	reg32 r1228 (rst, clk, in, r1228_out);
	reg32 r1229 (rst, clk, in, r1229_out);
	reg32 r1230 (rst, clk, in, r1230_out);
	reg32 r1231 (rst, clk, in, r1231_out);
	reg32 r1232 (rst, clk, in, r1232_out);
	reg32 r1233 (rst, clk, in, r1233_out);
	reg32 r1234 (rst, clk, in, r1234_out);
	reg32 r1235 (rst, clk, in, r1235_out);
	reg32 r1236 (rst, clk, in, r1236_out);
	reg32 r1237 (rst, clk, in, r1237_out);
	reg32 r1238 (rst, clk, in, r1238_out);
	reg32 r1239 (rst, clk, in, r1239_out);
	reg32 r1240 (rst, clk, in, r1240_out);
	reg32 r1241 (rst, clk, in, r1241_out);
	reg32 r1242 (rst, clk, in, r1242_out);
	reg32 r1243 (rst, clk, in, r1243_out);
	reg32 r1244 (rst, clk, in, r1244_out);
	reg32 r1245 (rst, clk, in, r1245_out);
	reg32 r1246 (rst, clk, in, r1246_out);
	reg32 r1247 (rst, clk, in, r1247_out);
	reg32 r1248 (rst, clk, in, r1248_out);
	reg32 r1249 (rst, clk, in, r1249_out);
	reg32 r1250 (rst, clk, in, r1250_out);
	reg32 r1251 (rst, clk, in, r1251_out);
	reg32 r1252 (rst, clk, in, r1252_out);
	reg32 r1253 (rst, clk, in, r1253_out);
	reg32 r1254 (rst, clk, in, r1254_out);
	reg32 r1255 (rst, clk, in, r1255_out);
	reg32 r1256 (rst, clk, in, r1256_out);
	reg32 r1257 (rst, clk, in, r1257_out);
	reg32 r1258 (rst, clk, in, r1258_out);
	reg32 r1259 (rst, clk, in, r1259_out);
	reg32 r1260 (rst, clk, in, r1260_out);
	reg32 r1261 (rst, clk, in, r1261_out);
	reg32 r1262 (rst, clk, in, r1262_out);
	reg32 r1263 (rst, clk, in, r1263_out);
	reg32 r1264 (rst, clk, in, r1264_out);
	reg32 r1265 (rst, clk, in, r1265_out);
	reg32 r1266 (rst, clk, in, r1266_out);
	reg32 r1267 (rst, clk, in, r1267_out);
	reg32 r1268 (rst, clk, in, r1268_out);
	reg32 r1269 (rst, clk, in, r1269_out);
	reg32 r1270 (rst, clk, in, r1270_out);
	reg32 r1271 (rst, clk, in, r1271_out);
	reg32 r1272 (rst, clk, in, r1272_out);
	reg32 r1273 (rst, clk, in, r1273_out);
	reg32 r1274 (rst, clk, in, r1274_out);
	reg32 r1275 (rst, clk, in, r1275_out);
	reg32 r1276 (rst, clk, in, r1276_out);
	reg32 r1277 (rst, clk, in, r1277_out);
	reg32 r1278 (rst, clk, in, r1278_out);
	reg32 r1279 (rst, clk, in, r1279_out);
	reg32 r1280 (rst, clk, in, r1280_out);
	reg32 r1281 (rst, clk, in, r1281_out);
	reg32 r1282 (rst, clk, in, r1282_out);
	reg32 r1283 (rst, clk, in, r1283_out);
	reg32 r1284 (rst, clk, in, r1284_out);
	reg32 r1285 (rst, clk, in, r1285_out);
	reg32 r1286 (rst, clk, in, r1286_out);
	reg32 r1287 (rst, clk, in, r1287_out);
	reg32 r1288 (rst, clk, in, r1288_out);
	reg32 r1289 (rst, clk, in, r1289_out);
	reg32 r1290 (rst, clk, in, r1290_out);
	reg32 r1291 (rst, clk, in, r1291_out);
	reg32 r1292 (rst, clk, in, r1292_out);
	reg32 r1293 (rst, clk, in, r1293_out);
	reg32 r1294 (rst, clk, in, r1294_out);
	reg32 r1295 (rst, clk, in, r1295_out);
	reg32 r1296 (rst, clk, in, r1296_out);
	reg32 r1297 (rst, clk, in, r1297_out);
	reg32 r1298 (rst, clk, in, r1298_out);
	reg32 r1299 (rst, clk, in, r1299_out);
	reg32 r1300 (rst, clk, in, r1300_out);
	reg32 r1301 (rst, clk, in, r1301_out);
	reg32 r1302 (rst, clk, in, r1302_out);
	reg32 r1303 (rst, clk, in, r1303_out);
	reg32 r1304 (rst, clk, in, r1304_out);
	reg32 r1305 (rst, clk, in, r1305_out);
	reg32 r1306 (rst, clk, in, r1306_out);
	reg32 r1307 (rst, clk, in, r1307_out);
	reg32 r1308 (rst, clk, in, r1308_out);
	reg32 r1309 (rst, clk, in, r1309_out);
	reg32 r1310 (rst, clk, in, r1310_out);
	reg32 r1311 (rst, clk, in, r1311_out);
	reg32 r1312 (rst, clk, in, r1312_out);
	reg32 r1313 (rst, clk, in, r1313_out);
	reg32 r1314 (rst, clk, in, r1314_out);
	reg32 r1315 (rst, clk, in, r1315_out);
	reg32 r1316 (rst, clk, in, r1316_out);
	reg32 r1317 (rst, clk, in, r1317_out);
	reg32 r1318 (rst, clk, in, r1318_out);
	reg32 r1319 (rst, clk, in, r1319_out);
	reg32 r1320 (rst, clk, in, r1320_out);
	reg32 r1321 (rst, clk, in, r1321_out);
	reg32 r1322 (rst, clk, in, r1322_out);
	reg32 r1323 (rst, clk, in, r1323_out);
	reg32 r1324 (rst, clk, in, r1324_out);
	reg32 r1325 (rst, clk, in, r1325_out);
	reg32 r1326 (rst, clk, in, r1326_out);
	reg32 r1327 (rst, clk, in, r1327_out);
	reg32 r1328 (rst, clk, in, r1328_out);
	reg32 r1329 (rst, clk, in, r1329_out);
	reg32 r1330 (rst, clk, in, r1330_out);
	reg32 r1331 (rst, clk, in, r1331_out);
	reg32 r1332 (rst, clk, in, r1332_out);
	reg32 r1333 (rst, clk, in, r1333_out);
	reg32 r1334 (rst, clk, in, r1334_out);
	reg32 r1335 (rst, clk, in, r1335_out);
	reg32 r1336 (rst, clk, in, r1336_out);
	reg32 r1337 (rst, clk, in, r1337_out);
	reg32 r1338 (rst, clk, in, r1338_out);
	reg32 r1339 (rst, clk, in, r1339_out);
	reg32 r1340 (rst, clk, in, r1340_out);
	reg32 r1341 (rst, clk, in, r1341_out);
	reg32 r1342 (rst, clk, in, r1342_out);
	reg32 r1343 (rst, clk, in, r1343_out);
	reg32 r1344 (rst, clk, in, r1344_out);
	reg32 r1345 (rst, clk, in, r1345_out);
	reg32 r1346 (rst, clk, in, r1346_out);
	reg32 r1347 (rst, clk, in, r1347_out);
	reg32 r1348 (rst, clk, in, r1348_out);
	reg32 r1349 (rst, clk, in, r1349_out);
	reg32 r1350 (rst, clk, in, r1350_out);
	reg32 r1351 (rst, clk, in, r1351_out);
	reg32 r1352 (rst, clk, in, r1352_out);
	reg32 r1353 (rst, clk, in, r1353_out);
	reg32 r1354 (rst, clk, in, r1354_out);
	reg32 r1355 (rst, clk, in, r1355_out);
	reg32 r1356 (rst, clk, in, r1356_out);
	reg32 r1357 (rst, clk, in, r1357_out);
	reg32 r1358 (rst, clk, in, r1358_out);
	reg32 r1359 (rst, clk, in, r1359_out);
	reg32 r1360 (rst, clk, in, r1360_out);
	reg32 r1361 (rst, clk, in, r1361_out);
	reg32 r1362 (rst, clk, in, r1362_out);
	reg32 r1363 (rst, clk, in, r1363_out);
	reg32 r1364 (rst, clk, in, r1364_out);
	reg32 r1365 (rst, clk, in, r1365_out);
	reg32 r1366 (rst, clk, in, r1366_out);
	reg32 r1367 (rst, clk, in, r1367_out);
	reg32 r1368 (rst, clk, in, r1368_out);
	reg32 r1369 (rst, clk, in, r1369_out);
	reg32 r1370 (rst, clk, in, r1370_out);
	reg32 r1371 (rst, clk, in, r1371_out);
	reg32 r1372 (rst, clk, in, r1372_out);
	reg32 r1373 (rst, clk, in, r1373_out);
	reg32 r1374 (rst, clk, in, r1374_out);
	reg32 r1375 (rst, clk, in, r1375_out);
	reg32 r1376 (rst, clk, in, r1376_out);
	reg32 r1377 (rst, clk, in, r1377_out);
	reg32 r1378 (rst, clk, in, r1378_out);
	reg32 r1379 (rst, clk, in, r1379_out);
	reg32 r1380 (rst, clk, in, r1380_out);
	reg32 r1381 (rst, clk, in, r1381_out);
	reg32 r1382 (rst, clk, in, r1382_out);
	reg32 r1383 (rst, clk, in, r1383_out);
	reg32 r1384 (rst, clk, in, r1384_out);
	reg32 r1385 (rst, clk, in, r1385_out);
	reg32 r1386 (rst, clk, in, r1386_out);
	reg32 r1387 (rst, clk, in, r1387_out);
	reg32 r1388 (rst, clk, in, r1388_out);
	reg32 r1389 (rst, clk, in, r1389_out);
	reg32 r1390 (rst, clk, in, r1390_out);
	reg32 r1391 (rst, clk, in, r1391_out);
	reg32 r1392 (rst, clk, in, r1392_out);
	reg32 r1393 (rst, clk, in, r1393_out);
	reg32 r1394 (rst, clk, in, r1394_out);
	reg32 r1395 (rst, clk, in, r1395_out);
	reg32 r1396 (rst, clk, in, r1396_out);
	reg32 r1397 (rst, clk, in, r1397_out);
	reg32 r1398 (rst, clk, in, r1398_out);
	reg32 r1399 (rst, clk, in, r1399_out);
	reg32 r1400 (rst, clk, in, r1400_out);
	reg32 r1401 (rst, clk, in, r1401_out);
	reg32 r1402 (rst, clk, in, r1402_out);
	reg32 r1403 (rst, clk, in, r1403_out);
	reg32 r1404 (rst, clk, in, r1404_out);
	reg32 r1405 (rst, clk, in, r1405_out);
	reg32 r1406 (rst, clk, in, r1406_out);
	reg32 r1407 (rst, clk, in, r1407_out);
	reg32 r1408 (rst, clk, in, r1408_out);
	reg32 r1409 (rst, clk, in, r1409_out);
	reg32 r1410 (rst, clk, in, r1410_out);
	reg32 r1411 (rst, clk, in, r1411_out);
	reg32 r1412 (rst, clk, in, r1412_out);
	reg32 r1413 (rst, clk, in, r1413_out);
	reg32 r1414 (rst, clk, in, r1414_out);
	reg32 r1415 (rst, clk, in, r1415_out);
	reg32 r1416 (rst, clk, in, r1416_out);
	reg32 r1417 (rst, clk, in, r1417_out);
	reg32 r1418 (rst, clk, in, r1418_out);
	reg32 r1419 (rst, clk, in, r1419_out);
	reg32 r1420 (rst, clk, in, r1420_out);
	reg32 r1421 (rst, clk, in, r1421_out);
	reg32 r1422 (rst, clk, in, r1422_out);
	reg32 r1423 (rst, clk, in, r1423_out);
	reg32 r1424 (rst, clk, in, r1424_out);
	reg32 r1425 (rst, clk, in, r1425_out);
	reg32 r1426 (rst, clk, in, r1426_out);
	reg32 r1427 (rst, clk, in, r1427_out);
	reg32 r1428 (rst, clk, in, r1428_out);
	reg32 r1429 (rst, clk, in, r1429_out);
	reg32 r1430 (rst, clk, in, r1430_out);
	reg32 r1431 (rst, clk, in, r1431_out);
	reg32 r1432 (rst, clk, in, r1432_out);
	reg32 r1433 (rst, clk, in, r1433_out);
	reg32 r1434 (rst, clk, in, r1434_out);
	reg32 r1435 (rst, clk, in, r1435_out);
	reg32 r1436 (rst, clk, in, r1436_out);
	reg32 r1437 (rst, clk, in, r1437_out);
	reg32 r1438 (rst, clk, in, r1438_out);
	reg32 r1439 (rst, clk, in, r1439_out);
	reg32 r1440 (rst, clk, in, r1440_out);
	reg32 r1441 (rst, clk, in, r1441_out);
	reg32 r1442 (rst, clk, in, r1442_out);
	reg32 r1443 (rst, clk, in, r1443_out);
	reg32 r1444 (rst, clk, in, r1444_out);
	reg32 r1445 (rst, clk, in, r1445_out);
	reg32 r1446 (rst, clk, in, r1446_out);
	reg32 r1447 (rst, clk, in, r1447_out);
	reg32 r1448 (rst, clk, in, r1448_out);
	reg32 r1449 (rst, clk, in, r1449_out);
	reg32 r1450 (rst, clk, in, r1450_out);
	reg32 r1451 (rst, clk, in, r1451_out);
	reg32 r1452 (rst, clk, in, r1452_out);
	reg32 r1453 (rst, clk, in, r1453_out);
	reg32 r1454 (rst, clk, in, r1454_out);
	reg32 r1455 (rst, clk, in, r1455_out);
	reg32 r1456 (rst, clk, in, r1456_out);
	reg32 r1457 (rst, clk, in, r1457_out);
	reg32 r1458 (rst, clk, in, r1458_out);
	reg32 r1459 (rst, clk, in, r1459_out);
	reg32 r1460 (rst, clk, in, r1460_out);
	reg32 r1461 (rst, clk, in, r1461_out);
	reg32 r1462 (rst, clk, in, r1462_out);
	reg32 r1463 (rst, clk, in, r1463_out);
	reg32 r1464 (rst, clk, in, r1464_out);
	reg32 r1465 (rst, clk, in, r1465_out);
	reg32 r1466 (rst, clk, in, r1466_out);
	reg32 r1467 (rst, clk, in, r1467_out);
	reg32 r1468 (rst, clk, in, r1468_out);
	reg32 r1469 (rst, clk, in, r1469_out);
	reg32 r1470 (rst, clk, in, r1470_out);
	reg32 r1471 (rst, clk, in, r1471_out);
	reg32 r1472 (rst, clk, in, r1472_out);
	reg32 r1473 (rst, clk, in, r1473_out);
	reg32 r1474 (rst, clk, in, r1474_out);
	reg32 r1475 (rst, clk, in, r1475_out);
	reg32 r1476 (rst, clk, in, r1476_out);
	reg32 r1477 (rst, clk, in, r1477_out);
	reg32 r1478 (rst, clk, in, r1478_out);
	reg32 r1479 (rst, clk, in, r1479_out);
	reg32 r1480 (rst, clk, in, r1480_out);
	reg32 r1481 (rst, clk, in, r1481_out);
	reg32 r1482 (rst, clk, in, r1482_out);
	reg32 r1483 (rst, clk, in, r1483_out);
	reg32 r1484 (rst, clk, in, r1484_out);
	reg32 r1485 (rst, clk, in, r1485_out);
	reg32 r1486 (rst, clk, in, r1486_out);
	reg32 r1487 (rst, clk, in, r1487_out);
	reg32 r1488 (rst, clk, in, r1488_out);
	reg32 r1489 (rst, clk, in, r1489_out);
	reg32 r1490 (rst, clk, in, r1490_out);
	reg32 r1491 (rst, clk, in, r1491_out);
	reg32 r1492 (rst, clk, in, r1492_out);
	reg32 r1493 (rst, clk, in, r1493_out);
	reg32 r1494 (rst, clk, in, r1494_out);
	reg32 r1495 (rst, clk, in, r1495_out);
	reg32 r1496 (rst, clk, in, r1496_out);
	reg32 r1497 (rst, clk, in, r1497_out);
	reg32 r1498 (rst, clk, in, r1498_out);
	reg32 r1499 (rst, clk, in, r1499_out);
	reg32 r1500 (rst, clk, in, r1500_out);
	reg32 r1501 (rst, clk, in, r1501_out);
	reg32 r1502 (rst, clk, in, r1502_out);
	reg32 r1503 (rst, clk, in, r1503_out);
	reg32 r1504 (rst, clk, in, r1504_out);
	reg32 r1505 (rst, clk, in, r1505_out);
	reg32 r1506 (rst, clk, in, r1506_out);
	reg32 r1507 (rst, clk, in, r1507_out);
	reg32 r1508 (rst, clk, in, r1508_out);
	reg32 r1509 (rst, clk, in, r1509_out);
	reg32 r1510 (rst, clk, in, r1510_out);
	reg32 r1511 (rst, clk, in, r1511_out);
	reg32 r1512 (rst, clk, in, r1512_out);
	reg32 r1513 (rst, clk, in, r1513_out);
	reg32 r1514 (rst, clk, in, r1514_out);
	reg32 r1515 (rst, clk, in, r1515_out);
	reg32 r1516 (rst, clk, in, r1516_out);
	reg32 r1517 (rst, clk, in, r1517_out);
	reg32 r1518 (rst, clk, in, r1518_out);
	reg32 r1519 (rst, clk, in, r1519_out);
	reg32 r1520 (rst, clk, in, r1520_out);
	reg32 r1521 (rst, clk, in, r1521_out);
	reg32 r1522 (rst, clk, in, r1522_out);
	reg32 r1523 (rst, clk, in, r1523_out);
	reg32 r1524 (rst, clk, in, r1524_out);
	reg32 r1525 (rst, clk, in, r1525_out);
	reg32 r1526 (rst, clk, in, r1526_out);
	reg32 r1527 (rst, clk, in, r1527_out);
	reg32 r1528 (rst, clk, in, r1528_out);
	reg32 r1529 (rst, clk, in, r1529_out);
	reg32 r1530 (rst, clk, in, r1530_out);
	reg32 r1531 (rst, clk, in, r1531_out);
	reg32 r1532 (rst, clk, in, r1532_out);
	reg32 r1533 (rst, clk, in, r1533_out);
	reg32 r1534 (rst, clk, in, r1534_out);
	reg32 r1535 (rst, clk, in, r1535_out);
	reg32 r1536 (rst, clk, in, r1536_out);
	reg32 r1537 (rst, clk, in, r1537_out);
	reg32 r1538 (rst, clk, in, r1538_out);
	reg32 r1539 (rst, clk, in, r1539_out);
	reg32 r1540 (rst, clk, in, r1540_out);
	reg32 r1541 (rst, clk, in, r1541_out);
	reg32 r1542 (rst, clk, in, r1542_out);
	reg32 r1543 (rst, clk, in, r1543_out);
	reg32 r1544 (rst, clk, in, r1544_out);
	reg32 r1545 (rst, clk, in, r1545_out);
	reg32 r1546 (rst, clk, in, r1546_out);
	reg32 r1547 (rst, clk, in, r1547_out);
	reg32 r1548 (rst, clk, in, r1548_out);
	reg32 r1549 (rst, clk, in, r1549_out);
	reg32 r1550 (rst, clk, in, r1550_out);
	reg32 r1551 (rst, clk, in, r1551_out);
	reg32 r1552 (rst, clk, in, r1552_out);
	reg32 r1553 (rst, clk, in, r1553_out);
	reg32 r1554 (rst, clk, in, r1554_out);
	reg32 r1555 (rst, clk, in, r1555_out);
	reg32 r1556 (rst, clk, in, r1556_out);
	reg32 r1557 (rst, clk, in, r1557_out);
	reg32 r1558 (rst, clk, in, r1558_out);
	reg32 r1559 (rst, clk, in, r1559_out);
	reg32 r1560 (rst, clk, in, r1560_out);
	reg32 r1561 (rst, clk, in, r1561_out);
	reg32 r1562 (rst, clk, in, r1562_out);
	reg32 r1563 (rst, clk, in, r1563_out);
	reg32 r1564 (rst, clk, in, r1564_out);
	reg32 r1565 (rst, clk, in, r1565_out);
	reg32 r1566 (rst, clk, in, r1566_out);
	reg32 r1567 (rst, clk, in, r1567_out);
	reg32 r1568 (rst, clk, in, r1568_out);
	reg32 r1569 (rst, clk, in, r1569_out);
	reg32 r1570 (rst, clk, in, r1570_out);
	reg32 r1571 (rst, clk, in, r1571_out);
	reg32 r1572 (rst, clk, in, r1572_out);
	reg32 r1573 (rst, clk, in, r1573_out);
	reg32 r1574 (rst, clk, in, r1574_out);
	reg32 r1575 (rst, clk, in, r1575_out);
	reg32 r1576 (rst, clk, in, r1576_out);
	reg32 r1577 (rst, clk, in, r1577_out);
	reg32 r1578 (rst, clk, in, r1578_out);
	reg32 r1579 (rst, clk, in, r1579_out);
	reg32 r1580 (rst, clk, in, r1580_out);
	reg32 r1581 (rst, clk, in, r1581_out);
	reg32 r1582 (rst, clk, in, r1582_out);
	reg32 r1583 (rst, clk, in, r1583_out);
	reg32 r1584 (rst, clk, in, r1584_out);
	reg32 r1585 (rst, clk, in, r1585_out);
	reg32 r1586 (rst, clk, in, r1586_out);
	reg32 r1587 (rst, clk, in, r1587_out);
	reg32 r1588 (rst, clk, in, r1588_out);
	reg32 r1589 (rst, clk, in, r1589_out);
	reg32 r1590 (rst, clk, in, r1590_out);
	reg32 r1591 (rst, clk, in, r1591_out);
	reg32 r1592 (rst, clk, in, r1592_out);
	reg32 r1593 (rst, clk, in, r1593_out);
	reg32 r1594 (rst, clk, in, r1594_out);
	reg32 r1595 (rst, clk, in, r1595_out);
	reg32 r1596 (rst, clk, in, r1596_out);
	reg32 r1597 (rst, clk, in, r1597_out);
	reg32 r1598 (rst, clk, in, r1598_out);
	reg32 r1599 (rst, clk, in, r1599_out);
	reg32 r1600 (rst, clk, in, r1600_out);
	reg32 r1601 (rst, clk, in, r1601_out);
	reg32 r1602 (rst, clk, in, r1602_out);
	reg32 r1603 (rst, clk, in, r1603_out);
	reg32 r1604 (rst, clk, in, r1604_out);
	reg32 r1605 (rst, clk, in, r1605_out);
	reg32 r1606 (rst, clk, in, r1606_out);
	reg32 r1607 (rst, clk, in, r1607_out);
	reg32 r1608 (rst, clk, in, r1608_out);
	reg32 r1609 (rst, clk, in, r1609_out);
	reg32 r1610 (rst, clk, in, r1610_out);
	reg32 r1611 (rst, clk, in, r1611_out);
	reg32 r1612 (rst, clk, in, r1612_out);
	reg32 r1613 (rst, clk, in, r1613_out);
	reg32 r1614 (rst, clk, in, r1614_out);
	reg32 r1615 (rst, clk, in, r1615_out);
	reg32 r1616 (rst, clk, in, r1616_out);
	reg32 r1617 (rst, clk, in, r1617_out);
	reg32 r1618 (rst, clk, in, r1618_out);
	reg32 r1619 (rst, clk, in, r1619_out);
	reg32 r1620 (rst, clk, in, r1620_out);
	reg32 r1621 (rst, clk, in, r1621_out);
	reg32 r1622 (rst, clk, in, r1622_out);
	reg32 r1623 (rst, clk, in, r1623_out);
	reg32 r1624 (rst, clk, in, r1624_out);
	reg32 r1625 (rst, clk, in, r1625_out);
	reg32 r1626 (rst, clk, in, r1626_out);
	reg32 r1627 (rst, clk, in, r1627_out);
	reg32 r1628 (rst, clk, in, r1628_out);
	reg32 r1629 (rst, clk, in, r1629_out);
	reg32 r1630 (rst, clk, in, r1630_out);
	reg32 r1631 (rst, clk, in, r1631_out);
	reg32 r1632 (rst, clk, in, r1632_out);
	reg32 r1633 (rst, clk, in, r1633_out);
	reg32 r1634 (rst, clk, in, r1634_out);
	reg32 r1635 (rst, clk, in, r1635_out);
	reg32 r1636 (rst, clk, in, r1636_out);
	reg32 r1637 (rst, clk, in, r1637_out);
	reg32 r1638 (rst, clk, in, r1638_out);
	reg32 r1639 (rst, clk, in, r1639_out);
	reg32 r1640 (rst, clk, in, r1640_out);
	reg32 r1641 (rst, clk, in, r1641_out);
	reg32 r1642 (rst, clk, in, r1642_out);
	reg32 r1643 (rst, clk, in, r1643_out);
	reg32 r1644 (rst, clk, in, r1644_out);
	reg32 r1645 (rst, clk, in, r1645_out);
	reg32 r1646 (rst, clk, in, r1646_out);
	reg32 r1647 (rst, clk, in, r1647_out);
	reg32 r1648 (rst, clk, in, r1648_out);
	reg32 r1649 (rst, clk, in, r1649_out);
	reg32 r1650 (rst, clk, in, r1650_out);
	reg32 r1651 (rst, clk, in, r1651_out);
	reg32 r1652 (rst, clk, in, r1652_out);
	reg32 r1653 (rst, clk, in, r1653_out);
	reg32 r1654 (rst, clk, in, r1654_out);
	reg32 r1655 (rst, clk, in, r1655_out);
	reg32 r1656 (rst, clk, in, r1656_out);
	reg32 r1657 (rst, clk, in, r1657_out);
	reg32 r1658 (rst, clk, in, r1658_out);
	reg32 r1659 (rst, clk, in, r1659_out);
	reg32 r1660 (rst, clk, in, r1660_out);
	reg32 r1661 (rst, clk, in, r1661_out);
	reg32 r1662 (rst, clk, in, r1662_out);
	reg32 r1663 (rst, clk, in, r1663_out);
	reg32 r1664 (rst, clk, in, r1664_out);
	reg32 r1665 (rst, clk, in, r1665_out);
	reg32 r1666 (rst, clk, in, r1666_out);
	reg32 r1667 (rst, clk, in, r1667_out);
	reg32 r1668 (rst, clk, in, r1668_out);
	reg32 r1669 (rst, clk, in, r1669_out);
	reg32 r1670 (rst, clk, in, r1670_out);
	reg32 r1671 (rst, clk, in, r1671_out);
	reg32 r1672 (rst, clk, in, r1672_out);
	reg32 r1673 (rst, clk, in, r1673_out);
	reg32 r1674 (rst, clk, in, r1674_out);
	reg32 r1675 (rst, clk, in, r1675_out);
	reg32 r1676 (rst, clk, in, r1676_out);
	reg32 r1677 (rst, clk, in, r1677_out);
	reg32 r1678 (rst, clk, in, r1678_out);
	reg32 r1679 (rst, clk, in, r1679_out);
	reg32 r1680 (rst, clk, in, r1680_out);
	reg32 r1681 (rst, clk, in, r1681_out);
	reg32 r1682 (rst, clk, in, r1682_out);
	reg32 r1683 (rst, clk, in, r1683_out);
	reg32 r1684 (rst, clk, in, r1684_out);
	reg32 r1685 (rst, clk, in, r1685_out);
	reg32 r1686 (rst, clk, in, r1686_out);
	reg32 r1687 (rst, clk, in, r1687_out);
	reg32 r1688 (rst, clk, in, r1688_out);
	reg32 r1689 (rst, clk, in, r1689_out);
	reg32 r1690 (rst, clk, in, r1690_out);
	reg32 r1691 (rst, clk, in, r1691_out);
	reg32 r1692 (rst, clk, in, r1692_out);
	reg32 r1693 (rst, clk, in, r1693_out);
	reg32 r1694 (rst, clk, in, r1694_out);
	reg32 r1695 (rst, clk, in, r1695_out);
	reg32 r1696 (rst, clk, in, r1696_out);
	reg32 r1697 (rst, clk, in, r1697_out);
	reg32 r1698 (rst, clk, in, r1698_out);
	reg32 r1699 (rst, clk, in, r1699_out);
	reg32 r1700 (rst, clk, in, r1700_out);
	reg32 r1701 (rst, clk, in, r1701_out);
	reg32 r1702 (rst, clk, in, r1702_out);
	reg32 r1703 (rst, clk, in, r1703_out);
	reg32 r1704 (rst, clk, in, r1704_out);
	reg32 r1705 (rst, clk, in, r1705_out);
	reg32 r1706 (rst, clk, in, r1706_out);
	reg32 r1707 (rst, clk, in, r1707_out);
	reg32 r1708 (rst, clk, in, r1708_out);
	reg32 r1709 (rst, clk, in, r1709_out);
	reg32 r1710 (rst, clk, in, r1710_out);
	reg32 r1711 (rst, clk, in, r1711_out);
	reg32 r1712 (rst, clk, in, r1712_out);
	reg32 r1713 (rst, clk, in, r1713_out);
	reg32 r1714 (rst, clk, in, r1714_out);
	reg32 r1715 (rst, clk, in, r1715_out);
	reg32 r1716 (rst, clk, in, r1716_out);
	reg32 r1717 (rst, clk, in, r1717_out);
	reg32 r1718 (rst, clk, in, r1718_out);
	reg32 r1719 (rst, clk, in, r1719_out);
	reg32 r1720 (rst, clk, in, r1720_out);
	reg32 r1721 (rst, clk, in, r1721_out);
	reg32 r1722 (rst, clk, in, r1722_out);
	reg32 r1723 (rst, clk, in, r1723_out);
	reg32 r1724 (rst, clk, in, r1724_out);
	reg32 r1725 (rst, clk, in, r1725_out);
	reg32 r1726 (rst, clk, in, r1726_out);
	reg32 r1727 (rst, clk, in, r1727_out);
	reg32 r1728 (rst, clk, in, r1728_out);
	reg32 r1729 (rst, clk, in, r1729_out);
	reg32 r1730 (rst, clk, in, r1730_out);
	reg32 r1731 (rst, clk, in, r1731_out);
	reg32 r1732 (rst, clk, in, r1732_out);
	reg32 r1733 (rst, clk, in, r1733_out);
	reg32 r1734 (rst, clk, in, r1734_out);
	reg32 r1735 (rst, clk, in, r1735_out);
	reg32 r1736 (rst, clk, in, r1736_out);
	reg32 r1737 (rst, clk, in, r1737_out);
	reg32 r1738 (rst, clk, in, r1738_out);
	reg32 r1739 (rst, clk, in, r1739_out);
	reg32 r1740 (rst, clk, in, r1740_out);
	reg32 r1741 (rst, clk, in, r1741_out);
	reg32 r1742 (rst, clk, in, r1742_out);
	reg32 r1743 (rst, clk, in, r1743_out);
	reg32 r1744 (rst, clk, in, r1744_out);
	reg32 r1745 (rst, clk, in, r1745_out);
	reg32 r1746 (rst, clk, in, r1746_out);
	reg32 r1747 (rst, clk, in, r1747_out);
	reg32 r1748 (rst, clk, in, r1748_out);
	reg32 r1749 (rst, clk, in, r1749_out);
	reg32 r1750 (rst, clk, in, r1750_out);
	reg32 r1751 (rst, clk, in, r1751_out);
	reg32 r1752 (rst, clk, in, r1752_out);
	reg32 r1753 (rst, clk, in, r1753_out);
	reg32 r1754 (rst, clk, in, r1754_out);
	reg32 r1755 (rst, clk, in, r1755_out);
	reg32 r1756 (rst, clk, in, r1756_out);
	reg32 r1757 (rst, clk, in, r1757_out);
	reg32 r1758 (rst, clk, in, r1758_out);
	reg32 r1759 (rst, clk, in, r1759_out);
	reg32 r1760 (rst, clk, in, r1760_out);
	reg32 r1761 (rst, clk, in, r1761_out);
	reg32 r1762 (rst, clk, in, r1762_out);
	reg32 r1763 (rst, clk, in, r1763_out);
	reg32 r1764 (rst, clk, in, r1764_out);
	reg32 r1765 (rst, clk, in, r1765_out);
	reg32 r1766 (rst, clk, in, r1766_out);
	reg32 r1767 (rst, clk, in, r1767_out);
	reg32 r1768 (rst, clk, in, r1768_out);
	reg32 r1769 (rst, clk, in, r1769_out);
	reg32 r1770 (rst, clk, in, r1770_out);
	reg32 r1771 (rst, clk, in, r1771_out);
	reg32 r1772 (rst, clk, in, r1772_out);
	reg32 r1773 (rst, clk, in, r1773_out);
	reg32 r1774 (rst, clk, in, r1774_out);
	reg32 r1775 (rst, clk, in, r1775_out);
	reg32 r1776 (rst, clk, in, r1776_out);
	reg32 r1777 (rst, clk, in, r1777_out);
	reg32 r1778 (rst, clk, in, r1778_out);
	reg32 r1779 (rst, clk, in, r1779_out);
	reg32 r1780 (rst, clk, in, r1780_out);
	reg32 r1781 (rst, clk, in, r1781_out);
	reg32 r1782 (rst, clk, in, r1782_out);
	reg32 r1783 (rst, clk, in, r1783_out);
	reg32 r1784 (rst, clk, in, r1784_out);
	reg32 r1785 (rst, clk, in, r1785_out);
	reg32 r1786 (rst, clk, in, r1786_out);
	reg32 r1787 (rst, clk, in, r1787_out);
	reg32 r1788 (rst, clk, in, r1788_out);
	reg32 r1789 (rst, clk, in, r1789_out);
	reg32 r1790 (rst, clk, in, r1790_out);
	reg32 r1791 (rst, clk, in, r1791_out);
	reg32 r1792 (rst, clk, in, r1792_out);
	reg32 r1793 (rst, clk, in, r1793_out);
	reg32 r1794 (rst, clk, in, r1794_out);
	reg32 r1795 (rst, clk, in, r1795_out);
	reg32 r1796 (rst, clk, in, r1796_out);
	reg32 r1797 (rst, clk, in, r1797_out);
	reg32 r1798 (rst, clk, in, r1798_out);
	reg32 r1799 (rst, clk, in, r1799_out);
	reg32 r1800 (rst, clk, in, r1800_out);
	reg32 r1801 (rst, clk, in, r1801_out);
	reg32 r1802 (rst, clk, in, r1802_out);
	reg32 r1803 (rst, clk, in, r1803_out);
	reg32 r1804 (rst, clk, in, r1804_out);
	reg32 r1805 (rst, clk, in, r1805_out);
	reg32 r1806 (rst, clk, in, r1806_out);
	reg32 r1807 (rst, clk, in, r1807_out);
	reg32 r1808 (rst, clk, in, r1808_out);
	reg32 r1809 (rst, clk, in, r1809_out);
	reg32 r1810 (rst, clk, in, r1810_out);
	reg32 r1811 (rst, clk, in, r1811_out);
	reg32 r1812 (rst, clk, in, r1812_out);
	reg32 r1813 (rst, clk, in, r1813_out);
	reg32 r1814 (rst, clk, in, r1814_out);
	reg32 r1815 (rst, clk, in, r1815_out);
	reg32 r1816 (rst, clk, in, r1816_out);
	reg32 r1817 (rst, clk, in, r1817_out);
	reg32 r1818 (rst, clk, in, r1818_out);
	reg32 r1819 (rst, clk, in, r1819_out);
	reg32 r1820 (rst, clk, in, r1820_out);
	reg32 r1821 (rst, clk, in, r1821_out);
	reg32 r1822 (rst, clk, in, r1822_out);
	reg32 r1823 (rst, clk, in, r1823_out);
	reg32 r1824 (rst, clk, in, r1824_out);
	reg32 r1825 (rst, clk, in, r1825_out);
	reg32 r1826 (rst, clk, in, r1826_out);
	reg32 r1827 (rst, clk, in, r1827_out);
	reg32 r1828 (rst, clk, in, r1828_out);
	reg32 r1829 (rst, clk, in, r1829_out);
	reg32 r1830 (rst, clk, in, r1830_out);
	reg32 r1831 (rst, clk, in, r1831_out);
	reg32 r1832 (rst, clk, in, r1832_out);
	reg32 r1833 (rst, clk, in, r1833_out);
	reg32 r1834 (rst, clk, in, r1834_out);
	reg32 r1835 (rst, clk, in, r1835_out);
	reg32 r1836 (rst, clk, in, r1836_out);
	reg32 r1837 (rst, clk, in, r1837_out);
	reg32 r1838 (rst, clk, in, r1838_out);
	reg32 r1839 (rst, clk, in, r1839_out);
	reg32 r1840 (rst, clk, in, r1840_out);
	reg32 r1841 (rst, clk, in, r1841_out);
	reg32 r1842 (rst, clk, in, r1842_out);
	reg32 r1843 (rst, clk, in, r1843_out);
	reg32 r1844 (rst, clk, in, r1844_out);
	reg32 r1845 (rst, clk, in, r1845_out);
	reg32 r1846 (rst, clk, in, r1846_out);
	reg32 r1847 (rst, clk, in, r1847_out);
	reg32 r1848 (rst, clk, in, r1848_out);
	reg32 r1849 (rst, clk, in, r1849_out);
	reg32 r1850 (rst, clk, in, r1850_out);
	reg32 r1851 (rst, clk, in, r1851_out);
	reg32 r1852 (rst, clk, in, r1852_out);
	reg32 r1853 (rst, clk, in, r1853_out);
	reg32 r1854 (rst, clk, in, r1854_out);
	reg32 r1855 (rst, clk, in, r1855_out);
	reg32 r1856 (rst, clk, in, r1856_out);
	reg32 r1857 (rst, clk, in, r1857_out);
	reg32 r1858 (rst, clk, in, r1858_out);
	reg32 r1859 (rst, clk, in, r1859_out);
	reg32 r1860 (rst, clk, in, r1860_out);
	reg32 r1861 (rst, clk, in, r1861_out);
	reg32 r1862 (rst, clk, in, r1862_out);
	reg32 r1863 (rst, clk, in, r1863_out);
	reg32 r1864 (rst, clk, in, r1864_out);
	reg32 r1865 (rst, clk, in, r1865_out);
	reg32 r1866 (rst, clk, in, r1866_out);
	reg32 r1867 (rst, clk, in, r1867_out);
	reg32 r1868 (rst, clk, in, r1868_out);
	reg32 r1869 (rst, clk, in, r1869_out);
	reg32 r1870 (rst, clk, in, r1870_out);
	reg32 r1871 (rst, clk, in, r1871_out);
	reg32 r1872 (rst, clk, in, r1872_out);
	reg32 r1873 (rst, clk, in, r1873_out);
	reg32 r1874 (rst, clk, in, r1874_out);
	reg32 r1875 (rst, clk, in, r1875_out);
	reg32 r1876 (rst, clk, in, r1876_out);
	reg32 r1877 (rst, clk, in, r1877_out);
	reg32 r1878 (rst, clk, in, r1878_out);
	reg32 r1879 (rst, clk, in, r1879_out);
	reg32 r1880 (rst, clk, in, r1880_out);
	reg32 r1881 (rst, clk, in, r1881_out);
	reg32 r1882 (rst, clk, in, r1882_out);
	reg32 r1883 (rst, clk, in, r1883_out);
	reg32 r1884 (rst, clk, in, r1884_out);
	reg32 r1885 (rst, clk, in, r1885_out);
	reg32 r1886 (rst, clk, in, r1886_out);
	reg32 r1887 (rst, clk, in, r1887_out);
	reg32 r1888 (rst, clk, in, r1888_out);
	reg32 r1889 (rst, clk, in, r1889_out);
	reg32 r1890 (rst, clk, in, r1890_out);
	reg32 r1891 (rst, clk, in, r1891_out);
	reg32 r1892 (rst, clk, in, r1892_out);
	reg32 r1893 (rst, clk, in, r1893_out);
	reg32 r1894 (rst, clk, in, r1894_out);
	reg32 r1895 (rst, clk, in, r1895_out);
	reg32 r1896 (rst, clk, in, r1896_out);
	reg32 r1897 (rst, clk, in, r1897_out);
	reg32 r1898 (rst, clk, in, r1898_out);
	reg32 r1899 (rst, clk, in, r1899_out);
	reg32 r1900 (rst, clk, in, r1900_out);
	reg32 r1901 (rst, clk, in, r1901_out);
	reg32 r1902 (rst, clk, in, r1902_out);
	reg32 r1903 (rst, clk, in, r1903_out);
	reg32 r1904 (rst, clk, in, r1904_out);
	reg32 r1905 (rst, clk, in, r1905_out);
	reg32 r1906 (rst, clk, in, r1906_out);
	reg32 r1907 (rst, clk, in, r1907_out);
	reg32 r1908 (rst, clk, in, r1908_out);
	reg32 r1909 (rst, clk, in, r1909_out);
	reg32 r1910 (rst, clk, in, r1910_out);
	reg32 r1911 (rst, clk, in, r1911_out);
	reg32 r1912 (rst, clk, in, r1912_out);
	reg32 r1913 (rst, clk, in, r1913_out);
	reg32 r1914 (rst, clk, in, r1914_out);
	reg32 r1915 (rst, clk, in, r1915_out);
	reg32 r1916 (rst, clk, in, r1916_out);
	reg32 r1917 (rst, clk, in, r1917_out);
	reg32 r1918 (rst, clk, in, r1918_out);
	reg32 r1919 (rst, clk, in, r1919_out);
	reg32 r1920 (rst, clk, in, r1920_out);
	reg32 r1921 (rst, clk, in, r1921_out);
	reg32 r1922 (rst, clk, in, r1922_out);
	reg32 r1923 (rst, clk, in, r1923_out);
	reg32 r1924 (rst, clk, in, r1924_out);
	reg32 r1925 (rst, clk, in, r1925_out);
	reg32 r1926 (rst, clk, in, r1926_out);
	reg32 r1927 (rst, clk, in, r1927_out);
	reg32 r1928 (rst, clk, in, r1928_out);
	reg32 r1929 (rst, clk, in, r1929_out);
	reg32 r1930 (rst, clk, in, r1930_out);
	reg32 r1931 (rst, clk, in, r1931_out);
	reg32 r1932 (rst, clk, in, r1932_out);
	reg32 r1933 (rst, clk, in, r1933_out);
	reg32 r1934 (rst, clk, in, r1934_out);
	reg32 r1935 (rst, clk, in, r1935_out);
	reg32 r1936 (rst, clk, in, r1936_out);
	reg32 r1937 (rst, clk, in, r1937_out);
	reg32 r1938 (rst, clk, in, r1938_out);
	reg32 r1939 (rst, clk, in, r1939_out);
	reg32 r1940 (rst, clk, in, r1940_out);
	reg32 r1941 (rst, clk, in, r1941_out);
	reg32 r1942 (rst, clk, in, r1942_out);
	reg32 r1943 (rst, clk, in, r1943_out);
	reg32 r1944 (rst, clk, in, r1944_out);
	reg32 r1945 (rst, clk, in, r1945_out);
	reg32 r1946 (rst, clk, in, r1946_out);
	reg32 r1947 (rst, clk, in, r1947_out);
	reg32 r1948 (rst, clk, in, r1948_out);
	reg32 r1949 (rst, clk, in, r1949_out);
	reg32 r1950 (rst, clk, in, r1950_out);
	reg32 r1951 (rst, clk, in, r1951_out);
	reg32 r1952 (rst, clk, in, r1952_out);
	reg32 r1953 (rst, clk, in, r1953_out);
	reg32 r1954 (rst, clk, in, r1954_out);
	reg32 r1955 (rst, clk, in, r1955_out);
	reg32 r1956 (rst, clk, in, r1956_out);
	reg32 r1957 (rst, clk, in, r1957_out);
	reg32 r1958 (rst, clk, in, r1958_out);
	reg32 r1959 (rst, clk, in, r1959_out);
	reg32 r1960 (rst, clk, in, r1960_out);
	reg32 r1961 (rst, clk, in, r1961_out);
	reg32 r1962 (rst, clk, in, r1962_out);
	reg32 r1963 (rst, clk, in, r1963_out);
	reg32 r1964 (rst, clk, in, r1964_out);
	reg32 r1965 (rst, clk, in, r1965_out);
	reg32 r1966 (rst, clk, in, r1966_out);
	reg32 r1967 (rst, clk, in, r1967_out);
	reg32 r1968 (rst, clk, in, r1968_out);
	reg32 r1969 (rst, clk, in, r1969_out);
	reg32 r1970 (rst, clk, in, r1970_out);
	reg32 r1971 (rst, clk, in, r1971_out);
	reg32 r1972 (rst, clk, in, r1972_out);
	reg32 r1973 (rst, clk, in, r1973_out);
	reg32 r1974 (rst, clk, in, r1974_out);
	reg32 r1975 (rst, clk, in, r1975_out);
	reg32 r1976 (rst, clk, in, r1976_out);
	reg32 r1977 (rst, clk, in, r1977_out);
	reg32 r1978 (rst, clk, in, r1978_out);
	reg32 r1979 (rst, clk, in, r1979_out);
	reg32 r1980 (rst, clk, in, r1980_out);
	reg32 r1981 (rst, clk, in, r1981_out);
	reg32 r1982 (rst, clk, in, r1982_out);
	reg32 r1983 (rst, clk, in, r1983_out);
	reg32 r1984 (rst, clk, in, r1984_out);
	reg32 r1985 (rst, clk, in, r1985_out);
	reg32 r1986 (rst, clk, in, r1986_out);
	reg32 r1987 (rst, clk, in, r1987_out);
	reg32 r1988 (rst, clk, in, r1988_out);
	reg32 r1989 (rst, clk, in, r1989_out);
	reg32 r1990 (rst, clk, in, r1990_out);
	reg32 r1991 (rst, clk, in, r1991_out);
	reg32 r1992 (rst, clk, in, r1992_out);
	reg32 r1993 (rst, clk, in, r1993_out);
	reg32 r1994 (rst, clk, in, r1994_out);
	reg32 r1995 (rst, clk, in, r1995_out);
	reg32 r1996 (rst, clk, in, r1996_out);
	reg32 r1997 (rst, clk, in, r1997_out);
	reg32 r1998 (rst, clk, in, r1998_out);
	reg32 r1999 (rst, clk, in, r1999_out);
	reg32 r2000 (rst, clk, in, r2000_out);
	reg32 r2001 (rst, clk, in, r2001_out);
	reg32 r2002 (rst, clk, in, r2002_out);
	reg32 r2003 (rst, clk, in, r2003_out);
	reg32 r2004 (rst, clk, in, r2004_out);
	reg32 r2005 (rst, clk, in, r2005_out);
	reg32 r2006 (rst, clk, in, r2006_out);
	reg32 r2007 (rst, clk, in, r2007_out);
	reg32 r2008 (rst, clk, in, r2008_out);
	reg32 r2009 (rst, clk, in, r2009_out);
	reg32 r2010 (rst, clk, in, r2010_out);
	reg32 r2011 (rst, clk, in, r2011_out);
	reg32 r2012 (rst, clk, in, r2012_out);
	reg32 r2013 (rst, clk, in, r2013_out);
	reg32 r2014 (rst, clk, in, r2014_out);
	reg32 r2015 (rst, clk, in, r2015_out);
	reg32 r2016 (rst, clk, in, r2016_out);
	reg32 r2017 (rst, clk, in, r2017_out);
	reg32 r2018 (rst, clk, in, r2018_out);
	reg32 r2019 (rst, clk, in, r2019_out);
	reg32 r2020 (rst, clk, in, r2020_out);
	reg32 r2021 (rst, clk, in, r2021_out);
	reg32 r2022 (rst, clk, in, r2022_out);
	reg32 r2023 (rst, clk, in, r2023_out);
	reg32 r2024 (rst, clk, in, r2024_out);
	reg32 r2025 (rst, clk, in, r2025_out);
	reg32 r2026 (rst, clk, in, r2026_out);
	reg32 r2027 (rst, clk, in, r2027_out);
	reg32 r2028 (rst, clk, in, r2028_out);
	reg32 r2029 (rst, clk, in, r2029_out);
	reg32 r2030 (rst, clk, in, r2030_out);
	reg32 r2031 (rst, clk, in, r2031_out);
	reg32 r2032 (rst, clk, in, r2032_out);
	reg32 r2033 (rst, clk, in, r2033_out);
	reg32 r2034 (rst, clk, in, r2034_out);
	reg32 r2035 (rst, clk, in, r2035_out);
	reg32 r2036 (rst, clk, in, r2036_out);
	reg32 r2037 (rst, clk, in, r2037_out);
	reg32 r2038 (rst, clk, in, r2038_out);
	reg32 r2039 (rst, clk, in, r2039_out);
	reg32 r2040 (rst, clk, in, r2040_out);
	reg32 r2041 (rst, clk, in, r2041_out);
	reg32 r2042 (rst, clk, in, r2042_out);
	reg32 r2043 (rst, clk, in, r2043_out);
	reg32 r2044 (rst, clk, in, r2044_out);
	reg32 r2045 (rst, clk, in, r2045_out);
	reg32 r2046 (rst, clk, in, r2046_out);
	reg32 r2047 (rst, clk, in, r2047_out);
	reg32 r2048 (rst, clk, in, r2048_out);
	reg32 r2049 (rst, clk, in, r2049_out);
	reg32 r2050 (rst, clk, in, r2050_out);
	reg32 r2051 (rst, clk, in, r2051_out);
	reg32 r2052 (rst, clk, in, r2052_out);
	reg32 r2053 (rst, clk, in, r2053_out);
	reg32 r2054 (rst, clk, in, r2054_out);
	reg32 r2055 (rst, clk, in, r2055_out);
	reg32 r2056 (rst, clk, in, r2056_out);
	reg32 r2057 (rst, clk, in, r2057_out);
	reg32 r2058 (rst, clk, in, r2058_out);
	reg32 r2059 (rst, clk, in, r2059_out);
	reg32 r2060 (rst, clk, in, r2060_out);
	reg32 r2061 (rst, clk, in, r2061_out);
	reg32 r2062 (rst, clk, in, r2062_out);
	reg32 r2063 (rst, clk, in, r2063_out);
	reg32 r2064 (rst, clk, in, r2064_out);
	reg32 r2065 (rst, clk, in, r2065_out);
	reg32 r2066 (rst, clk, in, r2066_out);
	reg32 r2067 (rst, clk, in, r2067_out);
	reg32 r2068 (rst, clk, in, r2068_out);
	reg32 r2069 (rst, clk, in, r2069_out);
	reg32 r2070 (rst, clk, in, r2070_out);
	reg32 r2071 (rst, clk, in, r2071_out);
	reg32 r2072 (rst, clk, in, r2072_out);
	reg32 r2073 (rst, clk, in, r2073_out);
	reg32 r2074 (rst, clk, in, r2074_out);
	reg32 r2075 (rst, clk, in, r2075_out);
	reg32 r2076 (rst, clk, in, r2076_out);
	reg32 r2077 (rst, clk, in, r2077_out);
	reg32 r2078 (rst, clk, in, r2078_out);
	reg32 r2079 (rst, clk, in, r2079_out);
	reg32 r2080 (rst, clk, in, r2080_out);
	reg32 r2081 (rst, clk, in, r2081_out);
	reg32 r2082 (rst, clk, in, r2082_out);
	reg32 r2083 (rst, clk, in, r2083_out);
	reg32 r2084 (rst, clk, in, r2084_out);
	reg32 r2085 (rst, clk, in, r2085_out);
	reg32 r2086 (rst, clk, in, r2086_out);
	reg32 r2087 (rst, clk, in, r2087_out);
	reg32 r2088 (rst, clk, in, r2088_out);
	reg32 r2089 (rst, clk, in, r2089_out);
	reg32 r2090 (rst, clk, in, r2090_out);
	reg32 r2091 (rst, clk, in, r2091_out);
	reg32 r2092 (rst, clk, in, r2092_out);
	reg32 r2093 (rst, clk, in, r2093_out);
	reg32 r2094 (rst, clk, in, r2094_out);
	reg32 r2095 (rst, clk, in, r2095_out);
	reg32 r2096 (rst, clk, in, r2096_out);
	reg32 r2097 (rst, clk, in, r2097_out);
	reg32 r2098 (rst, clk, in, r2098_out);
	reg32 r2099 (rst, clk, in, r2099_out);
	reg32 r2100 (rst, clk, in, r2100_out);
	reg32 r2101 (rst, clk, in, r2101_out);
	reg32 r2102 (rst, clk, in, r2102_out);
	reg32 r2103 (rst, clk, in, r2103_out);
	reg32 r2104 (rst, clk, in, r2104_out);
	reg32 r2105 (rst, clk, in, r2105_out);
	reg32 r2106 (rst, clk, in, r2106_out);
	reg32 r2107 (rst, clk, in, r2107_out);
	reg32 r2108 (rst, clk, in, r2108_out);
	reg32 r2109 (rst, clk, in, r2109_out);
	reg32 r2110 (rst, clk, in, r2110_out);
	reg32 r2111 (rst, clk, in, r2111_out);
	reg32 r2112 (rst, clk, in, r2112_out);
	reg32 r2113 (rst, clk, in, r2113_out);
	reg32 r2114 (rst, clk, in, r2114_out);
	reg32 r2115 (rst, clk, in, r2115_out);
	reg32 r2116 (rst, clk, in, r2116_out);
	reg32 r2117 (rst, clk, in, r2117_out);
	reg32 r2118 (rst, clk, in, r2118_out);
	reg32 r2119 (rst, clk, in, r2119_out);
	reg32 r2120 (rst, clk, in, r2120_out);
	reg32 r2121 (rst, clk, in, r2121_out);
	reg32 r2122 (rst, clk, in, r2122_out);
	reg32 r2123 (rst, clk, in, r2123_out);
	reg32 r2124 (rst, clk, in, r2124_out);
	reg32 r2125 (rst, clk, in, r2125_out);
	reg32 r2126 (rst, clk, in, r2126_out);
	reg32 r2127 (rst, clk, in, r2127_out);
	reg32 r2128 (rst, clk, in, r2128_out);
	reg32 r2129 (rst, clk, in, r2129_out);
	reg32 r2130 (rst, clk, in, r2130_out);
	reg32 r2131 (rst, clk, in, r2131_out);
	reg32 r2132 (rst, clk, in, r2132_out);
	reg32 r2133 (rst, clk, in, r2133_out);
	reg32 r2134 (rst, clk, in, r2134_out);
	reg32 r2135 (rst, clk, in, r2135_out);
	reg32 r2136 (rst, clk, in, r2136_out);
	reg32 r2137 (rst, clk, in, r2137_out);
	reg32 r2138 (rst, clk, in, r2138_out);
	reg32 r2139 (rst, clk, in, r2139_out);
	reg32 r2140 (rst, clk, in, r2140_out);
	reg32 r2141 (rst, clk, in, r2141_out);
	reg32 r2142 (rst, clk, in, r2142_out);
	reg32 r2143 (rst, clk, in, r2143_out);
	reg32 r2144 (rst, clk, in, r2144_out);
	reg32 r2145 (rst, clk, in, r2145_out);
	reg32 r2146 (rst, clk, in, r2146_out);
	reg32 r2147 (rst, clk, in, r2147_out);
	reg32 r2148 (rst, clk, in, r2148_out);
	reg32 r2149 (rst, clk, in, r2149_out);
	reg32 r2150 (rst, clk, in, r2150_out);
	reg32 r2151 (rst, clk, in, r2151_out);
	reg32 r2152 (rst, clk, in, r2152_out);
	reg32 r2153 (rst, clk, in, r2153_out);
	reg32 r2154 (rst, clk, in, r2154_out);
	reg32 r2155 (rst, clk, in, r2155_out);
	reg32 r2156 (rst, clk, in, r2156_out);
	reg32 r2157 (rst, clk, in, r2157_out);
	reg32 r2158 (rst, clk, in, r2158_out);
	reg32 r2159 (rst, clk, in, r2159_out);
	reg32 r2160 (rst, clk, in, r2160_out);
	reg32 r2161 (rst, clk, in, r2161_out);
	reg32 r2162 (rst, clk, in, r2162_out);
	reg32 r2163 (rst, clk, in, r2163_out);
	reg32 r2164 (rst, clk, in, r2164_out);
	reg32 r2165 (rst, clk, in, r2165_out);
	reg32 r2166 (rst, clk, in, r2166_out);
	reg32 r2167 (rst, clk, in, r2167_out);
	reg32 r2168 (rst, clk, in, r2168_out);
	reg32 r2169 (rst, clk, in, r2169_out);
	reg32 r2170 (rst, clk, in, r2170_out);
	reg32 r2171 (rst, clk, in, r2171_out);
	reg32 r2172 (rst, clk, in, r2172_out);
	reg32 r2173 (rst, clk, in, r2173_out);
	reg32 r2174 (rst, clk, in, r2174_out);
	reg32 r2175 (rst, clk, in, r2175_out);
	reg32 r2176 (rst, clk, in, r2176_out);
	reg32 r2177 (rst, clk, in, r2177_out);
	reg32 r2178 (rst, clk, in, r2178_out);
	reg32 r2179 (rst, clk, in, r2179_out);
	reg32 r2180 (rst, clk, in, r2180_out);
	reg32 r2181 (rst, clk, in, r2181_out);
	reg32 r2182 (rst, clk, in, r2182_out);
	reg32 r2183 (rst, clk, in, r2183_out);
	reg32 r2184 (rst, clk, in, r2184_out);
	reg32 r2185 (rst, clk, in, r2185_out);
	reg32 r2186 (rst, clk, in, r2186_out);
	reg32 r2187 (rst, clk, in, r2187_out);
	reg32 r2188 (rst, clk, in, r2188_out);
	reg32 r2189 (rst, clk, in, r2189_out);
	reg32 r2190 (rst, clk, in, r2190_out);
	reg32 r2191 (rst, clk, in, r2191_out);
	reg32 r2192 (rst, clk, in, r2192_out);
	reg32 r2193 (rst, clk, in, r2193_out);
	reg32 r2194 (rst, clk, in, r2194_out);
	reg32 r2195 (rst, clk, in, r2195_out);
	reg32 r2196 (rst, clk, in, r2196_out);
	reg32 r2197 (rst, clk, in, r2197_out);
	reg32 r2198 (rst, clk, in, r2198_out);
	reg32 r2199 (rst, clk, in, r2199_out);
	reg32 r2200 (rst, clk, in, r2200_out);
	reg32 r2201 (rst, clk, in, r2201_out);
	reg32 r2202 (rst, clk, in, r2202_out);
	reg32 r2203 (rst, clk, in, r2203_out);
	reg32 r2204 (rst, clk, in, r2204_out);
	reg32 r2205 (rst, clk, in, r2205_out);
	reg32 r2206 (rst, clk, in, r2206_out);
	reg32 r2207 (rst, clk, in, r2207_out);
	reg32 r2208 (rst, clk, in, r2208_out);
	reg32 r2209 (rst, clk, in, r2209_out);
	reg32 r2210 (rst, clk, in, r2210_out);
	reg32 r2211 (rst, clk, in, r2211_out);
	reg32 r2212 (rst, clk, in, r2212_out);
	reg32 r2213 (rst, clk, in, r2213_out);
	reg32 r2214 (rst, clk, in, r2214_out);
	reg32 r2215 (rst, clk, in, r2215_out);
	reg32 r2216 (rst, clk, in, r2216_out);
	reg32 r2217 (rst, clk, in, r2217_out);
	reg32 r2218 (rst, clk, in, r2218_out);
	reg32 r2219 (rst, clk, in, r2219_out);
	reg32 r2220 (rst, clk, in, r2220_out);
	reg32 r2221 (rst, clk, in, r2221_out);
	reg32 r2222 (rst, clk, in, r2222_out);
	reg32 r2223 (rst, clk, in, r2223_out);
	reg32 r2224 (rst, clk, in, r2224_out);
	reg32 r2225 (rst, clk, in, r2225_out);
	reg32 r2226 (rst, clk, in, r2226_out);
	reg32 r2227 (rst, clk, in, r2227_out);
	reg32 r2228 (rst, clk, in, r2228_out);
	reg32 r2229 (rst, clk, in, r2229_out);
	reg32 r2230 (rst, clk, in, r2230_out);
	reg32 r2231 (rst, clk, in, r2231_out);
	reg32 r2232 (rst, clk, in, r2232_out);
	reg32 r2233 (rst, clk, in, r2233_out);
	reg32 r2234 (rst, clk, in, r2234_out);
	reg32 r2235 (rst, clk, in, r2235_out);
	reg32 r2236 (rst, clk, in, r2236_out);
	reg32 r2237 (rst, clk, in, r2237_out);
	reg32 r2238 (rst, clk, in, r2238_out);
	reg32 r2239 (rst, clk, in, r2239_out);
	reg32 r2240 (rst, clk, in, r2240_out);
	reg32 r2241 (rst, clk, in, r2241_out);
	reg32 r2242 (rst, clk, in, r2242_out);
	reg32 r2243 (rst, clk, in, r2243_out);
	reg32 r2244 (rst, clk, in, r2244_out);
	reg32 r2245 (rst, clk, in, r2245_out);
	reg32 r2246 (rst, clk, in, r2246_out);
	reg32 r2247 (rst, clk, in, r2247_out);
	reg32 r2248 (rst, clk, in, r2248_out);
	reg32 r2249 (rst, clk, in, r2249_out);
	reg32 r2250 (rst, clk, in, r2250_out);
	reg32 r2251 (rst, clk, in, r2251_out);
	reg32 r2252 (rst, clk, in, r2252_out);
	reg32 r2253 (rst, clk, in, r2253_out);
	reg32 r2254 (rst, clk, in, r2254_out);
	reg32 r2255 (rst, clk, in, r2255_out);
	reg32 r2256 (rst, clk, in, r2256_out);
	reg32 r2257 (rst, clk, in, r2257_out);
	reg32 r2258 (rst, clk, in, r2258_out);
	reg32 r2259 (rst, clk, in, r2259_out);
	reg32 r2260 (rst, clk, in, r2260_out);
	reg32 r2261 (rst, clk, in, r2261_out);
	reg32 r2262 (rst, clk, in, r2262_out);
	reg32 r2263 (rst, clk, in, r2263_out);
	reg32 r2264 (rst, clk, in, r2264_out);
	reg32 r2265 (rst, clk, in, r2265_out);
	reg32 r2266 (rst, clk, in, r2266_out);
	reg32 r2267 (rst, clk, in, r2267_out);
	reg32 r2268 (rst, clk, in, r2268_out);
	reg32 r2269 (rst, clk, in, r2269_out);
	reg32 r2270 (rst, clk, in, r2270_out);
	reg32 r2271 (rst, clk, in, r2271_out);
	reg32 r2272 (rst, clk, in, r2272_out);
	reg32 r2273 (rst, clk, in, r2273_out);
	reg32 r2274 (rst, clk, in, r2274_out);
	reg32 r2275 (rst, clk, in, r2275_out);
	reg32 r2276 (rst, clk, in, r2276_out);
	reg32 r2277 (rst, clk, in, r2277_out);
	reg32 r2278 (rst, clk, in, r2278_out);
	reg32 r2279 (rst, clk, in, r2279_out);
	reg32 r2280 (rst, clk, in, r2280_out);
	reg32 r2281 (rst, clk, in, r2281_out);
	reg32 r2282 (rst, clk, in, r2282_out);
	reg32 r2283 (rst, clk, in, r2283_out);
	reg32 r2284 (rst, clk, in, r2284_out);
	reg32 r2285 (rst, clk, in, r2285_out);
	reg32 r2286 (rst, clk, in, r2286_out);
	reg32 r2287 (rst, clk, in, r2287_out);
	reg32 r2288 (rst, clk, in, r2288_out);
	reg32 r2289 (rst, clk, in, r2289_out);
	reg32 r2290 (rst, clk, in, r2290_out);
	reg32 r2291 (rst, clk, in, r2291_out);
	reg32 r2292 (rst, clk, in, r2292_out);
	reg32 r2293 (rst, clk, in, r2293_out);
	reg32 r2294 (rst, clk, in, r2294_out);
	reg32 r2295 (rst, clk, in, r2295_out);
	reg32 r2296 (rst, clk, in, r2296_out);
	reg32 r2297 (rst, clk, in, r2297_out);
	reg32 r2298 (rst, clk, in, r2298_out);
	reg32 r2299 (rst, clk, in, r2299_out);
	reg32 r2300 (rst, clk, in, r2300_out);
	reg32 r2301 (rst, clk, in, r2301_out);
	reg32 r2302 (rst, clk, in, r2302_out);
	reg32 r2303 (rst, clk, in, r2303_out);
	reg32 r2304 (rst, clk, in, r2304_out);
	reg32 r2305 (rst, clk, in, r2305_out);
	reg32 r2306 (rst, clk, in, r2306_out);
	reg32 r2307 (rst, clk, in, r2307_out);
	reg32 r2308 (rst, clk, in, r2308_out);
	reg32 r2309 (rst, clk, in, r2309_out);
	reg32 r2310 (rst, clk, in, r2310_out);
	reg32 r2311 (rst, clk, in, r2311_out);
	reg32 r2312 (rst, clk, in, r2312_out);
	reg32 r2313 (rst, clk, in, r2313_out);
	reg32 r2314 (rst, clk, in, r2314_out);
	reg32 r2315 (rst, clk, in, r2315_out);
	reg32 r2316 (rst, clk, in, r2316_out);
	reg32 r2317 (rst, clk, in, r2317_out);
	reg32 r2318 (rst, clk, in, r2318_out);
	reg32 r2319 (rst, clk, in, r2319_out);
	reg32 r2320 (rst, clk, in, r2320_out);
	reg32 r2321 (rst, clk, in, r2321_out);
	reg32 r2322 (rst, clk, in, r2322_out);
	reg32 r2323 (rst, clk, in, r2323_out);
	reg32 r2324 (rst, clk, in, r2324_out);
	reg32 r2325 (rst, clk, in, r2325_out);
	reg32 r2326 (rst, clk, in, r2326_out);
	reg32 r2327 (rst, clk, in, r2327_out);
	reg32 r2328 (rst, clk, in, r2328_out);
	reg32 r2329 (rst, clk, in, r2329_out);
	reg32 r2330 (rst, clk, in, r2330_out);
	reg32 r2331 (rst, clk, in, r2331_out);
	reg32 r2332 (rst, clk, in, r2332_out);
	reg32 r2333 (rst, clk, in, r2333_out);
	reg32 r2334 (rst, clk, in, r2334_out);
	reg32 r2335 (rst, clk, in, r2335_out);
	reg32 r2336 (rst, clk, in, r2336_out);
	reg32 r2337 (rst, clk, in, r2337_out);
	reg32 r2338 (rst, clk, in, r2338_out);
	reg32 r2339 (rst, clk, in, r2339_out);
	reg32 r2340 (rst, clk, in, r2340_out);
	reg32 r2341 (rst, clk, in, r2341_out);
	reg32 r2342 (rst, clk, in, r2342_out);
	reg32 r2343 (rst, clk, in, r2343_out);
	reg32 r2344 (rst, clk, in, r2344_out);
	reg32 r2345 (rst, clk, in, r2345_out);
	reg32 r2346 (rst, clk, in, r2346_out);
	reg32 r2347 (rst, clk, in, r2347_out);
	reg32 r2348 (rst, clk, in, r2348_out);
	reg32 r2349 (rst, clk, in, r2349_out);
	reg32 r2350 (rst, clk, in, r2350_out);
	reg32 r2351 (rst, clk, in, r2351_out);
	reg32 r2352 (rst, clk, in, r2352_out);
	reg32 r2353 (rst, clk, in, r2353_out);
	reg32 r2354 (rst, clk, in, r2354_out);
	reg32 r2355 (rst, clk, in, r2355_out);
	reg32 r2356 (rst, clk, in, r2356_out);
	reg32 r2357 (rst, clk, in, r2357_out);
	reg32 r2358 (rst, clk, in, r2358_out);
	reg32 r2359 (rst, clk, in, r2359_out);
	reg32 r2360 (rst, clk, in, r2360_out);
	reg32 r2361 (rst, clk, in, r2361_out);
	reg32 r2362 (rst, clk, in, r2362_out);
	reg32 r2363 (rst, clk, in, r2363_out);
	reg32 r2364 (rst, clk, in, r2364_out);
	reg32 r2365 (rst, clk, in, r2365_out);
	reg32 r2366 (rst, clk, in, r2366_out);
	reg32 r2367 (rst, clk, in, r2367_out);
	reg32 r2368 (rst, clk, in, r2368_out);
	reg32 r2369 (rst, clk, in, r2369_out);
	reg32 r2370 (rst, clk, in, r2370_out);
	reg32 r2371 (rst, clk, in, r2371_out);
	reg32 r2372 (rst, clk, in, r2372_out);
	reg32 r2373 (rst, clk, in, r2373_out);
	reg32 r2374 (rst, clk, in, r2374_out);
	reg32 r2375 (rst, clk, in, r2375_out);
	reg32 r2376 (rst, clk, in, r2376_out);
	reg32 r2377 (rst, clk, in, r2377_out);
	reg32 r2378 (rst, clk, in, r2378_out);
	reg32 r2379 (rst, clk, in, r2379_out);
	reg32 r2380 (rst, clk, in, r2380_out);
	reg32 r2381 (rst, clk, in, r2381_out);
	reg32 r2382 (rst, clk, in, r2382_out);
	reg32 r2383 (rst, clk, in, r2383_out);
	reg32 r2384 (rst, clk, in, r2384_out);
	reg32 r2385 (rst, clk, in, r2385_out);
	reg32 r2386 (rst, clk, in, r2386_out);
	reg32 r2387 (rst, clk, in, r2387_out);
	reg32 r2388 (rst, clk, in, r2388_out);
	reg32 r2389 (rst, clk, in, r2389_out);
	reg32 r2390 (rst, clk, in, r2390_out);
	reg32 r2391 (rst, clk, in, r2391_out);
	reg32 r2392 (rst, clk, in, r2392_out);
	reg32 r2393 (rst, clk, in, r2393_out);
	reg32 r2394 (rst, clk, in, r2394_out);
	reg32 r2395 (rst, clk, in, r2395_out);
	reg32 r2396 (rst, clk, in, r2396_out);
	reg32 r2397 (rst, clk, in, r2397_out);
	reg32 r2398 (rst, clk, in, r2398_out);
	reg32 r2399 (rst, clk, in, r2399_out);
	reg32 r2400 (rst, clk, in, r2400_out);
	reg32 r2401 (rst, clk, in, r2401_out);
	reg32 r2402 (rst, clk, in, r2402_out);
	reg32 r2403 (rst, clk, in, r2403_out);
	reg32 r2404 (rst, clk, in, r2404_out);
	reg32 r2405 (rst, clk, in, r2405_out);
	reg32 r2406 (rst, clk, in, r2406_out);
	reg32 r2407 (rst, clk, in, r2407_out);
	reg32 r2408 (rst, clk, in, r2408_out);
	reg32 r2409 (rst, clk, in, r2409_out);
	reg32 r2410 (rst, clk, in, r2410_out);
	reg32 r2411 (rst, clk, in, r2411_out);
	reg32 r2412 (rst, clk, in, r2412_out);
	reg32 r2413 (rst, clk, in, r2413_out);
	reg32 r2414 (rst, clk, in, r2414_out);
	reg32 r2415 (rst, clk, in, r2415_out);
	reg32 r2416 (rst, clk, in, r2416_out);
	reg32 r2417 (rst, clk, in, r2417_out);
	reg32 r2418 (rst, clk, in, r2418_out);
	reg32 r2419 (rst, clk, in, r2419_out);
	reg32 r2420 (rst, clk, in, r2420_out);
	reg32 r2421 (rst, clk, in, r2421_out);
	reg32 r2422 (rst, clk, in, r2422_out);
	reg32 r2423 (rst, clk, in, r2423_out);
	reg32 r2424 (rst, clk, in, r2424_out);
	reg32 r2425 (rst, clk, in, r2425_out);
	reg32 r2426 (rst, clk, in, r2426_out);
	reg32 r2427 (rst, clk, in, r2427_out);
	reg32 r2428 (rst, clk, in, r2428_out);
	reg32 r2429 (rst, clk, in, r2429_out);
	reg32 r2430 (rst, clk, in, r2430_out);
	reg32 r2431 (rst, clk, in, r2431_out);
	reg32 r2432 (rst, clk, in, r2432_out);
	reg32 r2433 (rst, clk, in, r2433_out);
	reg32 r2434 (rst, clk, in, r2434_out);
	reg32 r2435 (rst, clk, in, r2435_out);
	reg32 r2436 (rst, clk, in, r2436_out);
	reg32 r2437 (rst, clk, in, r2437_out);
	reg32 r2438 (rst, clk, in, r2438_out);
	reg32 r2439 (rst, clk, in, r2439_out);
	reg32 r2440 (rst, clk, in, r2440_out);
	reg32 r2441 (rst, clk, in, r2441_out);
	reg32 r2442 (rst, clk, in, r2442_out);
	reg32 r2443 (rst, clk, in, r2443_out);
	reg32 r2444 (rst, clk, in, r2444_out);
	reg32 r2445 (rst, clk, in, r2445_out);
	reg32 r2446 (rst, clk, in, r2446_out);
	reg32 r2447 (rst, clk, in, r2447_out);
	reg32 r2448 (rst, clk, in, r2448_out);
	reg32 r2449 (rst, clk, in, r2449_out);
	reg32 r2450 (rst, clk, in, r2450_out);
	reg32 r2451 (rst, clk, in, r2451_out);
	reg32 r2452 (rst, clk, in, r2452_out);
	reg32 r2453 (rst, clk, in, r2453_out);
	reg32 r2454 (rst, clk, in, r2454_out);
	reg32 r2455 (rst, clk, in, r2455_out);
	reg32 r2456 (rst, clk, in, r2456_out);
	reg32 r2457 (rst, clk, in, r2457_out);
	reg32 r2458 (rst, clk, in, r2458_out);
	reg32 r2459 (rst, clk, in, r2459_out);
	reg32 r2460 (rst, clk, in, r2460_out);
	reg32 r2461 (rst, clk, in, r2461_out);
	reg32 r2462 (rst, clk, in, r2462_out);
	reg32 r2463 (rst, clk, in, r2463_out);
	reg32 r2464 (rst, clk, in, r2464_out);
	reg32 r2465 (rst, clk, in, r2465_out);
	reg32 r2466 (rst, clk, in, r2466_out);
	reg32 r2467 (rst, clk, in, r2467_out);
	reg32 r2468 (rst, clk, in, r2468_out);
	reg32 r2469 (rst, clk, in, r2469_out);
	reg32 r2470 (rst, clk, in, r2470_out);
	reg32 r2471 (rst, clk, in, r2471_out);
	reg32 r2472 (rst, clk, in, r2472_out);
	reg32 r2473 (rst, clk, in, r2473_out);
	reg32 r2474 (rst, clk, in, r2474_out);
	reg32 r2475 (rst, clk, in, r2475_out);
	reg32 r2476 (rst, clk, in, r2476_out);
	reg32 r2477 (rst, clk, in, r2477_out);
	reg32 r2478 (rst, clk, in, r2478_out);
	reg32 r2479 (rst, clk, in, r2479_out);
	reg32 r2480 (rst, clk, in, r2480_out);
	reg32 r2481 (rst, clk, in, r2481_out);
	reg32 r2482 (rst, clk, in, r2482_out);
	reg32 r2483 (rst, clk, in, r2483_out);
	reg32 r2484 (rst, clk, in, r2484_out);
	reg32 r2485 (rst, clk, in, r2485_out);
	reg32 r2486 (rst, clk, in, r2486_out);
	reg32 r2487 (rst, clk, in, r2487_out);
	reg32 r2488 (rst, clk, in, r2488_out);
	reg32 r2489 (rst, clk, in, r2489_out);
	reg32 r2490 (rst, clk, in, r2490_out);
	reg32 r2491 (rst, clk, in, r2491_out);
	reg32 r2492 (rst, clk, in, r2492_out);
	reg32 r2493 (rst, clk, in, r2493_out);
	reg32 r2494 (rst, clk, in, r2494_out);
	reg32 r2495 (rst, clk, in, r2495_out);
	reg32 r2496 (rst, clk, in, r2496_out);
	reg32 r2497 (rst, clk, in, r2497_out);
	reg32 r2498 (rst, clk, in, r2498_out);
	reg32 r2499 (rst, clk, in, r2499_out);
	reg32 r2500 (rst, clk, in, r2500_out);
	reg32 r2501 (rst, clk, in, r2501_out);
	reg32 r2502 (rst, clk, in, r2502_out);
	reg32 r2503 (rst, clk, in, r2503_out);
	reg32 r2504 (rst, clk, in, r2504_out);
	reg32 r2505 (rst, clk, in, r2505_out);
	reg32 r2506 (rst, clk, in, r2506_out);
	reg32 r2507 (rst, clk, in, r2507_out);
	reg32 r2508 (rst, clk, in, r2508_out);
	reg32 r2509 (rst, clk, in, r2509_out);
	reg32 r2510 (rst, clk, in, r2510_out);
	reg32 r2511 (rst, clk, in, r2511_out);
	reg32 r2512 (rst, clk, in, r2512_out);
	reg32 r2513 (rst, clk, in, r2513_out);
	reg32 r2514 (rst, clk, in, r2514_out);
	reg32 r2515 (rst, clk, in, r2515_out);
	reg32 r2516 (rst, clk, in, r2516_out);
	reg32 r2517 (rst, clk, in, r2517_out);
	reg32 r2518 (rst, clk, in, r2518_out);
	reg32 r2519 (rst, clk, in, r2519_out);
	reg32 r2520 (rst, clk, in, r2520_out);
	reg32 r2521 (rst, clk, in, r2521_out);
	reg32 r2522 (rst, clk, in, r2522_out);
	reg32 r2523 (rst, clk, in, r2523_out);
	reg32 r2524 (rst, clk, in, r2524_out);
	reg32 r2525 (rst, clk, in, r2525_out);
	reg32 r2526 (rst, clk, in, r2526_out);
	reg32 r2527 (rst, clk, in, r2527_out);
	reg32 r2528 (rst, clk, in, r2528_out);
	reg32 r2529 (rst, clk, in, r2529_out);
	reg32 r2530 (rst, clk, in, r2530_out);
	reg32 r2531 (rst, clk, in, r2531_out);
	reg32 r2532 (rst, clk, in, r2532_out);
	reg32 r2533 (rst, clk, in, r2533_out);
	reg32 r2534 (rst, clk, in, r2534_out);
	reg32 r2535 (rst, clk, in, r2535_out);
	reg32 r2536 (rst, clk, in, r2536_out);
	reg32 r2537 (rst, clk, in, r2537_out);
	reg32 r2538 (rst, clk, in, r2538_out);
	reg32 r2539 (rst, clk, in, r2539_out);
	reg32 r2540 (rst, clk, in, r2540_out);
	reg32 r2541 (rst, clk, in, r2541_out);
	reg32 r2542 (rst, clk, in, r2542_out);
	reg32 r2543 (rst, clk, in, r2543_out);
	reg32 r2544 (rst, clk, in, r2544_out);
	reg32 r2545 (rst, clk, in, r2545_out);
	reg32 r2546 (rst, clk, in, r2546_out);
	reg32 r2547 (rst, clk, in, r2547_out);
	reg32 r2548 (rst, clk, in, r2548_out);
	reg32 r2549 (rst, clk, in, r2549_out);
	reg32 r2550 (rst, clk, in, r2550_out);
	reg32 r2551 (rst, clk, in, r2551_out);
	reg32 r2552 (rst, clk, in, r2552_out);
	reg32 r2553 (rst, clk, in, r2553_out);
	reg32 r2554 (rst, clk, in, r2554_out);
	reg32 r2555 (rst, clk, in, r2555_out);
	reg32 r2556 (rst, clk, in, r2556_out);
	reg32 r2557 (rst, clk, in, r2557_out);
	reg32 r2558 (rst, clk, in, r2558_out);
	reg32 r2559 (rst, clk, in, r2559_out);
	reg32 r2560 (rst, clk, in, r2560_out);
	reg32 r2561 (rst, clk, in, r2561_out);
	reg32 r2562 (rst, clk, in, r2562_out);
	reg32 r2563 (rst, clk, in, r2563_out);
	reg32 r2564 (rst, clk, in, r2564_out);
	reg32 r2565 (rst, clk, in, r2565_out);
	reg32 r2566 (rst, clk, in, r2566_out);
	reg32 r2567 (rst, clk, in, r2567_out);
	reg32 r2568 (rst, clk, in, r2568_out);
	reg32 r2569 (rst, clk, in, r2569_out);
	reg32 r2570 (rst, clk, in, r2570_out);
	reg32 r2571 (rst, clk, in, r2571_out);
	reg32 r2572 (rst, clk, in, r2572_out);
	reg32 r2573 (rst, clk, in, r2573_out);
	reg32 r2574 (rst, clk, in, r2574_out);
	reg32 r2575 (rst, clk, in, r2575_out);
	reg32 r2576 (rst, clk, in, r2576_out);
	reg32 r2577 (rst, clk, in, r2577_out);
	reg32 r2578 (rst, clk, in, r2578_out);
	reg32 r2579 (rst, clk, in, r2579_out);
	reg32 r2580 (rst, clk, in, r2580_out);
	reg32 r2581 (rst, clk, in, r2581_out);
	reg32 r2582 (rst, clk, in, r2582_out);
	reg32 r2583 (rst, clk, in, r2583_out);
	reg32 r2584 (rst, clk, in, r2584_out);
	reg32 r2585 (rst, clk, in, r2585_out);
	reg32 r2586 (rst, clk, in, r2586_out);
	reg32 r2587 (rst, clk, in, r2587_out);
	reg32 r2588 (rst, clk, in, r2588_out);
	reg32 r2589 (rst, clk, in, r2589_out);
	reg32 r2590 (rst, clk, in, r2590_out);
	reg32 r2591 (rst, clk, in, r2591_out);
	reg32 r2592 (rst, clk, in, r2592_out);
	reg32 r2593 (rst, clk, in, r2593_out);
	reg32 r2594 (rst, clk, in, r2594_out);
	reg32 r2595 (rst, clk, in, r2595_out);
	reg32 r2596 (rst, clk, in, r2596_out);
	reg32 r2597 (rst, clk, in, r2597_out);
	reg32 r2598 (rst, clk, in, r2598_out);
	reg32 r2599 (rst, clk, in, r2599_out);
	reg32 r2600 (rst, clk, in, r2600_out);
	reg32 r2601 (rst, clk, in, r2601_out);
	reg32 r2602 (rst, clk, in, r2602_out);
	reg32 r2603 (rst, clk, in, r2603_out);
	reg32 r2604 (rst, clk, in, r2604_out);
	reg32 r2605 (rst, clk, in, r2605_out);
	reg32 r2606 (rst, clk, in, r2606_out);
	reg32 r2607 (rst, clk, in, r2607_out);
	reg32 r2608 (rst, clk, in, r2608_out);
	reg32 r2609 (rst, clk, in, r2609_out);
	reg32 r2610 (rst, clk, in, r2610_out);
	reg32 r2611 (rst, clk, in, r2611_out);
	reg32 r2612 (rst, clk, in, r2612_out);
	reg32 r2613 (rst, clk, in, r2613_out);
	reg32 r2614 (rst, clk, in, r2614_out);
	reg32 r2615 (rst, clk, in, r2615_out);
	reg32 r2616 (rst, clk, in, r2616_out);
	reg32 r2617 (rst, clk, in, r2617_out);
	reg32 r2618 (rst, clk, in, r2618_out);
	reg32 r2619 (rst, clk, in, r2619_out);
	reg32 r2620 (rst, clk, in, r2620_out);
	reg32 r2621 (rst, clk, in, r2621_out);
	reg32 r2622 (rst, clk, in, r2622_out);
	reg32 r2623 (rst, clk, in, r2623_out);
	reg32 r2624 (rst, clk, in, r2624_out);
	reg32 r2625 (rst, clk, in, r2625_out);
	reg32 r2626 (rst, clk, in, r2626_out);
	reg32 r2627 (rst, clk, in, r2627_out);
	reg32 r2628 (rst, clk, in, r2628_out);
	reg32 r2629 (rst, clk, in, r2629_out);
	reg32 r2630 (rst, clk, in, r2630_out);
	reg32 r2631 (rst, clk, in, r2631_out);
	reg32 r2632 (rst, clk, in, r2632_out);
	reg32 r2633 (rst, clk, in, r2633_out);
	reg32 r2634 (rst, clk, in, r2634_out);
	reg32 r2635 (rst, clk, in, r2635_out);
	reg32 r2636 (rst, clk, in, r2636_out);
	reg32 r2637 (rst, clk, in, r2637_out);
	reg32 r2638 (rst, clk, in, r2638_out);
	reg32 r2639 (rst, clk, in, r2639_out);
	reg32 r2640 (rst, clk, in, r2640_out);
	reg32 r2641 (rst, clk, in, r2641_out);
	reg32 r2642 (rst, clk, in, r2642_out);
	reg32 r2643 (rst, clk, in, r2643_out);
	reg32 r2644 (rst, clk, in, r2644_out);
	reg32 r2645 (rst, clk, in, r2645_out);
	reg32 r2646 (rst, clk, in, r2646_out);
	reg32 r2647 (rst, clk, in, r2647_out);
	reg32 r2648 (rst, clk, in, r2648_out);
	reg32 r2649 (rst, clk, in, r2649_out);
	reg32 r2650 (rst, clk, in, r2650_out);
	reg32 r2651 (rst, clk, in, r2651_out);
	reg32 r2652 (rst, clk, in, r2652_out);
	reg32 r2653 (rst, clk, in, r2653_out);
	reg32 r2654 (rst, clk, in, r2654_out);
	reg32 r2655 (rst, clk, in, r2655_out);
	reg32 r2656 (rst, clk, in, r2656_out);
	reg32 r2657 (rst, clk, in, r2657_out);
	reg32 r2658 (rst, clk, in, r2658_out);
	reg32 r2659 (rst, clk, in, r2659_out);
	reg32 r2660 (rst, clk, in, r2660_out);
	reg32 r2661 (rst, clk, in, r2661_out);
	reg32 r2662 (rst, clk, in, r2662_out);
	reg32 r2663 (rst, clk, in, r2663_out);
	reg32 r2664 (rst, clk, in, r2664_out);
	reg32 r2665 (rst, clk, in, r2665_out);
	reg32 r2666 (rst, clk, in, r2666_out);
	reg32 r2667 (rst, clk, in, r2667_out);
	reg32 r2668 (rst, clk, in, r2668_out);
	reg32 r2669 (rst, clk, in, r2669_out);
	reg32 r2670 (rst, clk, in, r2670_out);
	reg32 r2671 (rst, clk, in, r2671_out);
	reg32 r2672 (rst, clk, in, r2672_out);
	reg32 r2673 (rst, clk, in, r2673_out);
	reg32 r2674 (rst, clk, in, r2674_out);
	reg32 r2675 (rst, clk, in, r2675_out);
	reg32 r2676 (rst, clk, in, r2676_out);
	reg32 r2677 (rst, clk, in, r2677_out);
	reg32 r2678 (rst, clk, in, r2678_out);
	reg32 r2679 (rst, clk, in, r2679_out);
	reg32 r2680 (rst, clk, in, r2680_out);
	reg32 r2681 (rst, clk, in, r2681_out);
	reg32 r2682 (rst, clk, in, r2682_out);
	reg32 r2683 (rst, clk, in, r2683_out);
	reg32 r2684 (rst, clk, in, r2684_out);
	reg32 r2685 (rst, clk, in, r2685_out);
	reg32 r2686 (rst, clk, in, r2686_out);
	reg32 r2687 (rst, clk, in, r2687_out);
	reg32 r2688 (rst, clk, in, r2688_out);
	reg32 r2689 (rst, clk, in, r2689_out);
	reg32 r2690 (rst, clk, in, r2690_out);
	reg32 r2691 (rst, clk, in, r2691_out);
	reg32 r2692 (rst, clk, in, r2692_out);
	reg32 r2693 (rst, clk, in, r2693_out);
	reg32 r2694 (rst, clk, in, r2694_out);
	reg32 r2695 (rst, clk, in, r2695_out);
	reg32 r2696 (rst, clk, in, r2696_out);
	reg32 r2697 (rst, clk, in, r2697_out);
	reg32 r2698 (rst, clk, in, r2698_out);
	reg32 r2699 (rst, clk, in, r2699_out);
	reg32 r2700 (rst, clk, in, r2700_out);
	reg32 r2701 (rst, clk, in, r2701_out);
	reg32 r2702 (rst, clk, in, r2702_out);
	reg32 r2703 (rst, clk, in, r2703_out);
	reg32 r2704 (rst, clk, in, r2704_out);
	reg32 r2705 (rst, clk, in, r2705_out);
	reg32 r2706 (rst, clk, in, r2706_out);
	reg32 r2707 (rst, clk, in, r2707_out);
	reg32 r2708 (rst, clk, in, r2708_out);
	reg32 r2709 (rst, clk, in, r2709_out);
	reg32 r2710 (rst, clk, in, r2710_out);
	reg32 r2711 (rst, clk, in, r2711_out);
	reg32 r2712 (rst, clk, in, r2712_out);
	reg32 r2713 (rst, clk, in, r2713_out);
	reg32 r2714 (rst, clk, in, r2714_out);
	reg32 r2715 (rst, clk, in, r2715_out);
	reg32 r2716 (rst, clk, in, r2716_out);
	reg32 r2717 (rst, clk, in, r2717_out);
	reg32 r2718 (rst, clk, in, r2718_out);
	reg32 r2719 (rst, clk, in, r2719_out);
	reg32 r2720 (rst, clk, in, r2720_out);
	reg32 r2721 (rst, clk, in, r2721_out);
	reg32 r2722 (rst, clk, in, r2722_out);
	reg32 r2723 (rst, clk, in, r2723_out);
	reg32 r2724 (rst, clk, in, r2724_out);
	reg32 r2725 (rst, clk, in, r2725_out);
	reg32 r2726 (rst, clk, in, r2726_out);
	reg32 r2727 (rst, clk, in, r2727_out);
	reg32 r2728 (rst, clk, in, r2728_out);
	reg32 r2729 (rst, clk, in, r2729_out);
	reg32 r2730 (rst, clk, in, r2730_out);
	reg32 r2731 (rst, clk, in, r2731_out);
	reg32 r2732 (rst, clk, in, r2732_out);
	reg32 r2733 (rst, clk, in, r2733_out);
	reg32 r2734 (rst, clk, in, r2734_out);
	reg32 r2735 (rst, clk, in, r2735_out);
	reg32 r2736 (rst, clk, in, r2736_out);
	reg32 r2737 (rst, clk, in, r2737_out);
	reg32 r2738 (rst, clk, in, r2738_out);
	reg32 r2739 (rst, clk, in, r2739_out);
	reg32 r2740 (rst, clk, in, r2740_out);
	reg32 r2741 (rst, clk, in, r2741_out);
	reg32 r2742 (rst, clk, in, r2742_out);
	reg32 r2743 (rst, clk, in, r2743_out);
	reg32 r2744 (rst, clk, in, r2744_out);
	reg32 r2745 (rst, clk, in, r2745_out);
	reg32 r2746 (rst, clk, in, r2746_out);
	reg32 r2747 (rst, clk, in, r2747_out);
	reg32 r2748 (rst, clk, in, r2748_out);
	reg32 r2749 (rst, clk, in, r2749_out);
	reg32 r2750 (rst, clk, in, r2750_out);
	reg32 r2751 (rst, clk, in, r2751_out);
	reg32 r2752 (rst, clk, in, r2752_out);
	reg32 r2753 (rst, clk, in, r2753_out);
	reg32 r2754 (rst, clk, in, r2754_out);
	reg32 r2755 (rst, clk, in, r2755_out);
	reg32 r2756 (rst, clk, in, r2756_out);
	reg32 r2757 (rst, clk, in, r2757_out);
	reg32 r2758 (rst, clk, in, r2758_out);
	reg32 r2759 (rst, clk, in, r2759_out);
	reg32 r2760 (rst, clk, in, r2760_out);
	reg32 r2761 (rst, clk, in, r2761_out);
	reg32 r2762 (rst, clk, in, r2762_out);
	reg32 r2763 (rst, clk, in, r2763_out);
	reg32 r2764 (rst, clk, in, r2764_out);
	reg32 r2765 (rst, clk, in, r2765_out);
	reg32 r2766 (rst, clk, in, r2766_out);
	reg32 r2767 (rst, clk, in, r2767_out);
	reg32 r2768 (rst, clk, in, r2768_out);
	reg32 r2769 (rst, clk, in, r2769_out);
	reg32 r2770 (rst, clk, in, r2770_out);
	reg32 r2771 (rst, clk, in, r2771_out);
	reg32 r2772 (rst, clk, in, r2772_out);
	reg32 r2773 (rst, clk, in, r2773_out);
	reg32 r2774 (rst, clk, in, r2774_out);
	reg32 r2775 (rst, clk, in, r2775_out);
	reg32 r2776 (rst, clk, in, r2776_out);
	reg32 r2777 (rst, clk, in, r2777_out);
	reg32 r2778 (rst, clk, in, r2778_out);
	reg32 r2779 (rst, clk, in, r2779_out);
	reg32 r2780 (rst, clk, in, r2780_out);
	reg32 r2781 (rst, clk, in, r2781_out);
	reg32 r2782 (rst, clk, in, r2782_out);
	reg32 r2783 (rst, clk, in, r2783_out);
	reg32 r2784 (rst, clk, in, r2784_out);
	reg32 r2785 (rst, clk, in, r2785_out);
	reg32 r2786 (rst, clk, in, r2786_out);
	reg32 r2787 (rst, clk, in, r2787_out);
	reg32 r2788 (rst, clk, in, r2788_out);
	reg32 r2789 (rst, clk, in, r2789_out);
	reg32 r2790 (rst, clk, in, r2790_out);
	reg32 r2791 (rst, clk, in, r2791_out);
	reg32 r2792 (rst, clk, in, r2792_out);
	reg32 r2793 (rst, clk, in, r2793_out);
	reg32 r2794 (rst, clk, in, r2794_out);
	reg32 r2795 (rst, clk, in, r2795_out);
	reg32 r2796 (rst, clk, in, r2796_out);
	reg32 r2797 (rst, clk, in, r2797_out);
	reg32 r2798 (rst, clk, in, r2798_out);
	reg32 r2799 (rst, clk, in, r2799_out);
	reg32 r2800 (rst, clk, in, r2800_out);
	reg32 r2801 (rst, clk, in, r2801_out);
	reg32 r2802 (rst, clk, in, r2802_out);
	reg32 r2803 (rst, clk, in, r2803_out);
	reg32 r2804 (rst, clk, in, r2804_out);
	reg32 r2805 (rst, clk, in, r2805_out);
	reg32 r2806 (rst, clk, in, r2806_out);
	reg32 r2807 (rst, clk, in, r2807_out);
	reg32 r2808 (rst, clk, in, r2808_out);
	reg32 r2809 (rst, clk, in, r2809_out);
	reg32 r2810 (rst, clk, in, r2810_out);
	reg32 r2811 (rst, clk, in, r2811_out);
	reg32 r2812 (rst, clk, in, r2812_out);
	reg32 r2813 (rst, clk, in, r2813_out);
	reg32 r2814 (rst, clk, in, r2814_out);
	reg32 r2815 (rst, clk, in, r2815_out);
	reg32 r2816 (rst, clk, in, r2816_out);
	reg32 r2817 (rst, clk, in, r2817_out);
	reg32 r2818 (rst, clk, in, r2818_out);
	reg32 r2819 (rst, clk, in, r2819_out);
	reg32 r2820 (rst, clk, in, r2820_out);
	reg32 r2821 (rst, clk, in, r2821_out);
	reg32 r2822 (rst, clk, in, r2822_out);
	reg32 r2823 (rst, clk, in, r2823_out);
	reg32 r2824 (rst, clk, in, r2824_out);
	reg32 r2825 (rst, clk, in, r2825_out);
	reg32 r2826 (rst, clk, in, r2826_out);
	reg32 r2827 (rst, clk, in, r2827_out);
	reg32 r2828 (rst, clk, in, r2828_out);
	reg32 r2829 (rst, clk, in, r2829_out);
	reg32 r2830 (rst, clk, in, r2830_out);
	reg32 r2831 (rst, clk, in, r2831_out);
	reg32 r2832 (rst, clk, in, r2832_out);
	reg32 r2833 (rst, clk, in, r2833_out);
	reg32 r2834 (rst, clk, in, r2834_out);
	reg32 r2835 (rst, clk, in, r2835_out);
	reg32 r2836 (rst, clk, in, r2836_out);
	reg32 r2837 (rst, clk, in, r2837_out);
	reg32 r2838 (rst, clk, in, r2838_out);
	reg32 r2839 (rst, clk, in, r2839_out);
	reg32 r2840 (rst, clk, in, r2840_out);
	reg32 r2841 (rst, clk, in, r2841_out);
	reg32 r2842 (rst, clk, in, r2842_out);
	reg32 r2843 (rst, clk, in, r2843_out);
	reg32 r2844 (rst, clk, in, r2844_out);
	reg32 r2845 (rst, clk, in, r2845_out);
	reg32 r2846 (rst, clk, in, r2846_out);
	reg32 r2847 (rst, clk, in, r2847_out);
	reg32 r2848 (rst, clk, in, r2848_out);
	reg32 r2849 (rst, clk, in, r2849_out);
	reg32 r2850 (rst, clk, in, r2850_out);
	reg32 r2851 (rst, clk, in, r2851_out);
	reg32 r2852 (rst, clk, in, r2852_out);
	reg32 r2853 (rst, clk, in, r2853_out);
	reg32 r2854 (rst, clk, in, r2854_out);
	reg32 r2855 (rst, clk, in, r2855_out);
	reg32 r2856 (rst, clk, in, r2856_out);
	reg32 r2857 (rst, clk, in, r2857_out);
	reg32 r2858 (rst, clk, in, r2858_out);
	reg32 r2859 (rst, clk, in, r2859_out);
	reg32 r2860 (rst, clk, in, r2860_out);
	reg32 r2861 (rst, clk, in, r2861_out);
	reg32 r2862 (rst, clk, in, r2862_out);
	reg32 r2863 (rst, clk, in, r2863_out);
	reg32 r2864 (rst, clk, in, r2864_out);
	reg32 r2865 (rst, clk, in, r2865_out);
	reg32 r2866 (rst, clk, in, r2866_out);
	reg32 r2867 (rst, clk, in, r2867_out);
	reg32 r2868 (rst, clk, in, r2868_out);
	reg32 r2869 (rst, clk, in, r2869_out);
	reg32 r2870 (rst, clk, in, r2870_out);
	reg32 r2871 (rst, clk, in, r2871_out);
	reg32 r2872 (rst, clk, in, r2872_out);
	reg32 r2873 (rst, clk, in, r2873_out);
	reg32 r2874 (rst, clk, in, r2874_out);
	reg32 r2875 (rst, clk, in, r2875_out);
	reg32 r2876 (rst, clk, in, r2876_out);
	reg32 r2877 (rst, clk, in, r2877_out);
	reg32 r2878 (rst, clk, in, r2878_out);
	reg32 r2879 (rst, clk, in, r2879_out);
	reg32 r2880 (rst, clk, in, r2880_out);
	reg32 r2881 (rst, clk, in, r2881_out);
	reg32 r2882 (rst, clk, in, r2882_out);
	reg32 r2883 (rst, clk, in, r2883_out);
	reg32 r2884 (rst, clk, in, r2884_out);
	reg32 r2885 (rst, clk, in, r2885_out);
	reg32 r2886 (rst, clk, in, r2886_out);
	reg32 r2887 (rst, clk, in, r2887_out);
	reg32 r2888 (rst, clk, in, r2888_out);
	reg32 r2889 (rst, clk, in, r2889_out);
	reg32 r2890 (rst, clk, in, r2890_out);
	reg32 r2891 (rst, clk, in, r2891_out);
	reg32 r2892 (rst, clk, in, r2892_out);
	reg32 r2893 (rst, clk, in, r2893_out);
	reg32 r2894 (rst, clk, in, r2894_out);
	reg32 r2895 (rst, clk, in, r2895_out);
	reg32 r2896 (rst, clk, in, r2896_out);
	reg32 r2897 (rst, clk, in, r2897_out);
	reg32 r2898 (rst, clk, in, r2898_out);
	reg32 r2899 (rst, clk, in, r2899_out);
	reg32 r2900 (rst, clk, in, r2900_out);
	reg32 r2901 (rst, clk, in, r2901_out);
	reg32 r2902 (rst, clk, in, r2902_out);
	reg32 r2903 (rst, clk, in, r2903_out);
	reg32 r2904 (rst, clk, in, r2904_out);
	reg32 r2905 (rst, clk, in, r2905_out);
	reg32 r2906 (rst, clk, in, r2906_out);
	reg32 r2907 (rst, clk, in, r2907_out);
	reg32 r2908 (rst, clk, in, r2908_out);
	reg32 r2909 (rst, clk, in, r2909_out);
	reg32 r2910 (rst, clk, in, r2910_out);
	reg32 r2911 (rst, clk, in, r2911_out);
	reg32 r2912 (rst, clk, in, r2912_out);
	reg32 r2913 (rst, clk, in, r2913_out);
	reg32 r2914 (rst, clk, in, r2914_out);
	reg32 r2915 (rst, clk, in, r2915_out);
	reg32 r2916 (rst, clk, in, r2916_out);
	reg32 r2917 (rst, clk, in, r2917_out);
	reg32 r2918 (rst, clk, in, r2918_out);
	reg32 r2919 (rst, clk, in, r2919_out);
	reg32 r2920 (rst, clk, in, r2920_out);
	reg32 r2921 (rst, clk, in, r2921_out);
	reg32 r2922 (rst, clk, in, r2922_out);
	reg32 r2923 (rst, clk, in, r2923_out);
	reg32 r2924 (rst, clk, in, r2924_out);
	reg32 r2925 (rst, clk, in, r2925_out);
	reg32 r2926 (rst, clk, in, r2926_out);
	reg32 r2927 (rst, clk, in, r2927_out);
	reg32 r2928 (rst, clk, in, r2928_out);
	reg32 r2929 (rst, clk, in, r2929_out);
	reg32 r2930 (rst, clk, in, r2930_out);
	reg32 r2931 (rst, clk, in, r2931_out);
	reg32 r2932 (rst, clk, in, r2932_out);
	reg32 r2933 (rst, clk, in, r2933_out);
	reg32 r2934 (rst, clk, in, r2934_out);
	reg32 r2935 (rst, clk, in, r2935_out);
	reg32 r2936 (rst, clk, in, r2936_out);
	reg32 r2937 (rst, clk, in, r2937_out);
	reg32 r2938 (rst, clk, in, r2938_out);
	reg32 r2939 (rst, clk, in, r2939_out);
	reg32 r2940 (rst, clk, in, r2940_out);
	reg32 r2941 (rst, clk, in, r2941_out);
	reg32 r2942 (rst, clk, in, r2942_out);
	reg32 r2943 (rst, clk, in, r2943_out);
	reg32 r2944 (rst, clk, in, r2944_out);
	reg32 r2945 (rst, clk, in, r2945_out);
	reg32 r2946 (rst, clk, in, r2946_out);
	reg32 r2947 (rst, clk, in, r2947_out);
	reg32 r2948 (rst, clk, in, r2948_out);
	reg32 r2949 (rst, clk, in, r2949_out);
	reg32 r2950 (rst, clk, in, r2950_out);
	reg32 r2951 (rst, clk, in, r2951_out);
	reg32 r2952 (rst, clk, in, r2952_out);
	reg32 r2953 (rst, clk, in, r2953_out);
	reg32 r2954 (rst, clk, in, r2954_out);
	reg32 r2955 (rst, clk, in, r2955_out);
	reg32 r2956 (rst, clk, in, r2956_out);
	reg32 r2957 (rst, clk, in, r2957_out);
	reg32 r2958 (rst, clk, in, r2958_out);
	reg32 r2959 (rst, clk, in, r2959_out);
	reg32 r2960 (rst, clk, in, r2960_out);
	reg32 r2961 (rst, clk, in, r2961_out);
	reg32 r2962 (rst, clk, in, r2962_out);
	reg32 r2963 (rst, clk, in, r2963_out);
	reg32 r2964 (rst, clk, in, r2964_out);
	reg32 r2965 (rst, clk, in, r2965_out);
	reg32 r2966 (rst, clk, in, r2966_out);
	reg32 r2967 (rst, clk, in, r2967_out);
	reg32 r2968 (rst, clk, in, r2968_out);
	reg32 r2969 (rst, clk, in, r2969_out);
	reg32 r2970 (rst, clk, in, r2970_out);
	reg32 r2971 (rst, clk, in, r2971_out);
	reg32 r2972 (rst, clk, in, r2972_out);
	reg32 r2973 (rst, clk, in, r2973_out);
	reg32 r2974 (rst, clk, in, r2974_out);
	reg32 r2975 (rst, clk, in, r2975_out);
	reg32 r2976 (rst, clk, in, r2976_out);
	reg32 r2977 (rst, clk, in, r2977_out);
	reg32 r2978 (rst, clk, in, r2978_out);
	reg32 r2979 (rst, clk, in, r2979_out);
	reg32 r2980 (rst, clk, in, r2980_out);
	reg32 r2981 (rst, clk, in, r2981_out);
	reg32 r2982 (rst, clk, in, r2982_out);
	reg32 r2983 (rst, clk, in, r2983_out);
	reg32 r2984 (rst, clk, in, r2984_out);
	reg32 r2985 (rst, clk, in, r2985_out);
	reg32 r2986 (rst, clk, in, r2986_out);
	reg32 r2987 (rst, clk, in, r2987_out);
	reg32 r2988 (rst, clk, in, r2988_out);
	reg32 r2989 (rst, clk, in, r2989_out);
	reg32 r2990 (rst, clk, in, r2990_out);
	reg32 r2991 (rst, clk, in, r2991_out);
	reg32 r2992 (rst, clk, in, r2992_out);
	reg32 r2993 (rst, clk, in, r2993_out);
	reg32 r2994 (rst, clk, in, r2994_out);
	reg32 r2995 (rst, clk, in, r2995_out);
	reg32 r2996 (rst, clk, in, r2996_out);
	reg32 r2997 (rst, clk, in, r2997_out);
	reg32 r2998 (rst, clk, in, r2998_out);
	reg32 r2999 (rst, clk, in, r2999_out);
	reg32 r3000 (rst, clk, in, r3000_out);
	reg32 r3001 (rst, clk, in, r3001_out);
	reg32 r3002 (rst, clk, in, r3002_out);
	reg32 r3003 (rst, clk, in, r3003_out);
	reg32 r3004 (rst, clk, in, r3004_out);
	reg32 r3005 (rst, clk, in, r3005_out);
	reg32 r3006 (rst, clk, in, r3006_out);
	reg32 r3007 (rst, clk, in, r3007_out);
	reg32 r3008 (rst, clk, in, r3008_out);
	reg32 r3009 (rst, clk, in, r3009_out);
	reg32 r3010 (rst, clk, in, r3010_out);
	reg32 r3011 (rst, clk, in, r3011_out);
	reg32 r3012 (rst, clk, in, r3012_out);
	reg32 r3013 (rst, clk, in, r3013_out);
	reg32 r3014 (rst, clk, in, r3014_out);
	reg32 r3015 (rst, clk, in, r3015_out);
	reg32 r3016 (rst, clk, in, r3016_out);
	reg32 r3017 (rst, clk, in, r3017_out);
	reg32 r3018 (rst, clk, in, r3018_out);
	reg32 r3019 (rst, clk, in, r3019_out);
	reg32 r3020 (rst, clk, in, r3020_out);
	reg32 r3021 (rst, clk, in, r3021_out);
	reg32 r3022 (rst, clk, in, r3022_out);
	reg32 r3023 (rst, clk, in, r3023_out);
	reg32 r3024 (rst, clk, in, r3024_out);
	reg32 r3025 (rst, clk, in, r3025_out);
	reg32 r3026 (rst, clk, in, r3026_out);
	reg32 r3027 (rst, clk, in, r3027_out);
	reg32 r3028 (rst, clk, in, r3028_out);
	reg32 r3029 (rst, clk, in, r3029_out);
	reg32 r3030 (rst, clk, in, r3030_out);
	reg32 r3031 (rst, clk, in, r3031_out);
	reg32 r3032 (rst, clk, in, r3032_out);
	reg32 r3033 (rst, clk, in, r3033_out);
	reg32 r3034 (rst, clk, in, r3034_out);
	reg32 r3035 (rst, clk, in, r3035_out);
	reg32 r3036 (rst, clk, in, r3036_out);
	reg32 r3037 (rst, clk, in, r3037_out);
	reg32 r3038 (rst, clk, in, r3038_out);
	reg32 r3039 (rst, clk, in, r3039_out);
	reg32 r3040 (rst, clk, in, r3040_out);
	reg32 r3041 (rst, clk, in, r3041_out);
	reg32 r3042 (rst, clk, in, r3042_out);
	reg32 r3043 (rst, clk, in, r3043_out);
	reg32 r3044 (rst, clk, in, r3044_out);
	reg32 r3045 (rst, clk, in, r3045_out);
	reg32 r3046 (rst, clk, in, r3046_out);
	reg32 r3047 (rst, clk, in, r3047_out);
	reg32 r3048 (rst, clk, in, r3048_out);
	reg32 r3049 (rst, clk, in, r3049_out);
	reg32 r3050 (rst, clk, in, r3050_out);
	reg32 r3051 (rst, clk, in, r3051_out);
	reg32 r3052 (rst, clk, in, r3052_out);
	reg32 r3053 (rst, clk, in, r3053_out);
	reg32 r3054 (rst, clk, in, r3054_out);
	reg32 r3055 (rst, clk, in, r3055_out);
	reg32 r3056 (rst, clk, in, r3056_out);
	reg32 r3057 (rst, clk, in, r3057_out);
	reg32 r3058 (rst, clk, in, r3058_out);
	reg32 r3059 (rst, clk, in, r3059_out);
	reg32 r3060 (rst, clk, in, r3060_out);
	reg32 r3061 (rst, clk, in, r3061_out);
	reg32 r3062 (rst, clk, in, r3062_out);
	reg32 r3063 (rst, clk, in, r3063_out);
	reg32 r3064 (rst, clk, in, r3064_out);
	reg32 r3065 (rst, clk, in, r3065_out);
	reg32 r3066 (rst, clk, in, r3066_out);
	reg32 r3067 (rst, clk, in, r3067_out);
	reg32 r3068 (rst, clk, in, r3068_out);
	reg32 r3069 (rst, clk, in, r3069_out);
	reg32 r3070 (rst, clk, in, r3070_out);
	reg32 r3071 (rst, clk, in, r3071_out);
	reg32 r3072 (rst, clk, in, r3072_out);
	reg32 r3073 (rst, clk, in, r3073_out);
	reg32 r3074 (rst, clk, in, r3074_out);
	reg32 r3075 (rst, clk, in, r3075_out);
	reg32 r3076 (rst, clk, in, r3076_out);
	reg32 r3077 (rst, clk, in, r3077_out);
	reg32 r3078 (rst, clk, in, r3078_out);
	reg32 r3079 (rst, clk, in, r3079_out);
	reg32 r3080 (rst, clk, in, r3080_out);
	reg32 r3081 (rst, clk, in, r3081_out);
	reg32 r3082 (rst, clk, in, r3082_out);
	reg32 r3083 (rst, clk, in, r3083_out);
	reg32 r3084 (rst, clk, in, r3084_out);
	reg32 r3085 (rst, clk, in, r3085_out);
	reg32 r3086 (rst, clk, in, r3086_out);
	reg32 r3087 (rst, clk, in, r3087_out);
	reg32 r3088 (rst, clk, in, r3088_out);
	reg32 r3089 (rst, clk, in, r3089_out);
	reg32 r3090 (rst, clk, in, r3090_out);
	reg32 r3091 (rst, clk, in, r3091_out);
	reg32 r3092 (rst, clk, in, r3092_out);
	reg32 r3093 (rst, clk, in, r3093_out);
	reg32 r3094 (rst, clk, in, r3094_out);
	reg32 r3095 (rst, clk, in, r3095_out);
	reg32 r3096 (rst, clk, in, r3096_out);
	reg32 r3097 (rst, clk, in, r3097_out);
	reg32 r3098 (rst, clk, in, r3098_out);
	reg32 r3099 (rst, clk, in, r3099_out);
	reg32 r3100 (rst, clk, in, r3100_out);
	reg32 r3101 (rst, clk, in, r3101_out);
	reg32 r3102 (rst, clk, in, r3102_out);
	reg32 r3103 (rst, clk, in, r3103_out);
	reg32 r3104 (rst, clk, in, r3104_out);
	reg32 r3105 (rst, clk, in, r3105_out);
	reg32 r3106 (rst, clk, in, r3106_out);
	reg32 r3107 (rst, clk, in, r3107_out);
	reg32 r3108 (rst, clk, in, r3108_out);
	reg32 r3109 (rst, clk, in, r3109_out);
	reg32 r3110 (rst, clk, in, r3110_out);
	reg32 r3111 (rst, clk, in, r3111_out);
	reg32 r3112 (rst, clk, in, r3112_out);
	reg32 r3113 (rst, clk, in, r3113_out);
	reg32 r3114 (rst, clk, in, r3114_out);
	reg32 r3115 (rst, clk, in, r3115_out);
	reg32 r3116 (rst, clk, in, r3116_out);
	reg32 r3117 (rst, clk, in, r3117_out);
	reg32 r3118 (rst, clk, in, r3118_out);
	reg32 r3119 (rst, clk, in, r3119_out);
	reg32 r3120 (rst, clk, in, r3120_out);
	reg32 r3121 (rst, clk, in, r3121_out);
	reg32 r3122 (rst, clk, in, r3122_out);
	reg32 r3123 (rst, clk, in, r3123_out);
	reg32 r3124 (rst, clk, in, r3124_out);
	reg32 r3125 (rst, clk, in, r3125_out);
	reg32 r3126 (rst, clk, in, r3126_out);
	reg32 r3127 (rst, clk, in, r3127_out);
	reg32 r3128 (rst, clk, in, r3128_out);
	reg32 r3129 (rst, clk, in, r3129_out);
	reg32 r3130 (rst, clk, in, r3130_out);
	reg32 r3131 (rst, clk, in, r3131_out);
	reg32 r3132 (rst, clk, in, r3132_out);
	reg32 r3133 (rst, clk, in, r3133_out);
	reg32 r3134 (rst, clk, in, r3134_out);
	reg32 r3135 (rst, clk, in, r3135_out);
	reg32 r3136 (rst, clk, in, r3136_out);
	reg32 r3137 (rst, clk, in, r3137_out);
	reg32 r3138 (rst, clk, in, r3138_out);
	reg32 r3139 (rst, clk, in, r3139_out);
	reg32 r3140 (rst, clk, in, r3140_out);
	reg32 r3141 (rst, clk, in, r3141_out);
	reg32 r3142 (rst, clk, in, r3142_out);
	reg32 r3143 (rst, clk, in, r3143_out);
	reg32 r3144 (rst, clk, in, r3144_out);
	reg32 r3145 (rst, clk, in, r3145_out);
	reg32 r3146 (rst, clk, in, r3146_out);
	reg32 r3147 (rst, clk, in, r3147_out);
	reg32 r3148 (rst, clk, in, r3148_out);
	reg32 r3149 (rst, clk, in, r3149_out);
	reg32 r3150 (rst, clk, in, r3150_out);
	reg32 r3151 (rst, clk, in, r3151_out);
	reg32 r3152 (rst, clk, in, r3152_out);
	reg32 r3153 (rst, clk, in, r3153_out);
	reg32 r3154 (rst, clk, in, r3154_out);
	reg32 r3155 (rst, clk, in, r3155_out);
	reg32 r3156 (rst, clk, in, r3156_out);
	reg32 r3157 (rst, clk, in, r3157_out);
	reg32 r3158 (rst, clk, in, r3158_out);
	reg32 r3159 (rst, clk, in, r3159_out);
	reg32 r3160 (rst, clk, in, r3160_out);
	reg32 r3161 (rst, clk, in, r3161_out);
	reg32 r3162 (rst, clk, in, r3162_out);
	reg32 r3163 (rst, clk, in, r3163_out);
	reg32 r3164 (rst, clk, in, r3164_out);
	reg32 r3165 (rst, clk, in, r3165_out);
	reg32 r3166 (rst, clk, in, r3166_out);
	reg32 r3167 (rst, clk, in, r3167_out);
	reg32 r3168 (rst, clk, in, r3168_out);
	reg32 r3169 (rst, clk, in, r3169_out);
	reg32 r3170 (rst, clk, in, r3170_out);
	reg32 r3171 (rst, clk, in, r3171_out);
	reg32 r3172 (rst, clk, in, r3172_out);
	reg32 r3173 (rst, clk, in, r3173_out);
	reg32 r3174 (rst, clk, in, r3174_out);
	reg32 r3175 (rst, clk, in, r3175_out);
	reg32 r3176 (rst, clk, in, r3176_out);
	reg32 r3177 (rst, clk, in, r3177_out);
	reg32 r3178 (rst, clk, in, r3178_out);
	reg32 r3179 (rst, clk, in, r3179_out);
	reg32 r3180 (rst, clk, in, r3180_out);
	reg32 r3181 (rst, clk, in, r3181_out);
	reg32 r3182 (rst, clk, in, r3182_out);
	reg32 r3183 (rst, clk, in, r3183_out);
	reg32 r3184 (rst, clk, in, r3184_out);
	reg32 r3185 (rst, clk, in, r3185_out);
	reg32 r3186 (rst, clk, in, r3186_out);
	reg32 r3187 (rst, clk, in, r3187_out);
	reg32 r3188 (rst, clk, in, r3188_out);
	reg32 r3189 (rst, clk, in, r3189_out);
	reg32 r3190 (rst, clk, in, r3190_out);
	reg32 r3191 (rst, clk, in, r3191_out);
	reg32 r3192 (rst, clk, in, r3192_out);
	reg32 r3193 (rst, clk, in, r3193_out);
	reg32 r3194 (rst, clk, in, r3194_out);
	reg32 r3195 (rst, clk, in, r3195_out);
	reg32 r3196 (rst, clk, in, r3196_out);
	reg32 r3197 (rst, clk, in, r3197_out);
	reg32 r3198 (rst, clk, in, r3198_out);
	reg32 r3199 (rst, clk, in, r3199_out);
	reg32 r3200 (rst, clk, in, r3200_out);
	reg32 r3201 (rst, clk, in, r3201_out);
	reg32 r3202 (rst, clk, in, r3202_out);
	reg32 r3203 (rst, clk, in, r3203_out);
	reg32 r3204 (rst, clk, in, r3204_out);
	reg32 r3205 (rst, clk, in, r3205_out);
	reg32 r3206 (rst, clk, in, r3206_out);
	reg32 r3207 (rst, clk, in, r3207_out);
	reg32 r3208 (rst, clk, in, r3208_out);
	reg32 r3209 (rst, clk, in, r3209_out);
	reg32 r3210 (rst, clk, in, r3210_out);
	reg32 r3211 (rst, clk, in, r3211_out);
	reg32 r3212 (rst, clk, in, r3212_out);
	reg32 r3213 (rst, clk, in, r3213_out);
	reg32 r3214 (rst, clk, in, r3214_out);
	reg32 r3215 (rst, clk, in, r3215_out);
	reg32 r3216 (rst, clk, in, r3216_out);
	reg32 r3217 (rst, clk, in, r3217_out);
	reg32 r3218 (rst, clk, in, r3218_out);
	reg32 r3219 (rst, clk, in, r3219_out);
	reg32 r3220 (rst, clk, in, r3220_out);
	reg32 r3221 (rst, clk, in, r3221_out);
	reg32 r3222 (rst, clk, in, r3222_out);
	reg32 r3223 (rst, clk, in, r3223_out);
	reg32 r3224 (rst, clk, in, r3224_out);
	reg32 r3225 (rst, clk, in, r3225_out);
	reg32 r3226 (rst, clk, in, r3226_out);
	reg32 r3227 (rst, clk, in, r3227_out);
	reg32 r3228 (rst, clk, in, r3228_out);
	reg32 r3229 (rst, clk, in, r3229_out);
	reg32 r3230 (rst, clk, in, r3230_out);
	reg32 r3231 (rst, clk, in, r3231_out);
	reg32 r3232 (rst, clk, in, r3232_out);
	reg32 r3233 (rst, clk, in, r3233_out);
	reg32 r3234 (rst, clk, in, r3234_out);
	reg32 r3235 (rst, clk, in, r3235_out);
	reg32 r3236 (rst, clk, in, r3236_out);
	reg32 r3237 (rst, clk, in, r3237_out);
	reg32 r3238 (rst, clk, in, r3238_out);
	reg32 r3239 (rst, clk, in, r3239_out);
	reg32 r3240 (rst, clk, in, r3240_out);
	reg32 r3241 (rst, clk, in, r3241_out);
	reg32 r3242 (rst, clk, in, r3242_out);
	reg32 r3243 (rst, clk, in, r3243_out);
	reg32 r3244 (rst, clk, in, r3244_out);
	reg32 r3245 (rst, clk, in, r3245_out);
	reg32 r3246 (rst, clk, in, r3246_out);
	reg32 r3247 (rst, clk, in, r3247_out);
	reg32 r3248 (rst, clk, in, r3248_out);
	reg32 r3249 (rst, clk, in, r3249_out);
	reg32 r3250 (rst, clk, in, r3250_out);
	reg32 r3251 (rst, clk, in, r3251_out);
	reg32 r3252 (rst, clk, in, r3252_out);
	reg32 r3253 (rst, clk, in, r3253_out);
	reg32 r3254 (rst, clk, in, r3254_out);
	reg32 r3255 (rst, clk, in, r3255_out);
	reg32 r3256 (rst, clk, in, r3256_out);
	reg32 r3257 (rst, clk, in, r3257_out);
	reg32 r3258 (rst, clk, in, r3258_out);
	reg32 r3259 (rst, clk, in, r3259_out);
	reg32 r3260 (rst, clk, in, r3260_out);
	reg32 r3261 (rst, clk, in, r3261_out);
	reg32 r3262 (rst, clk, in, r3262_out);
	reg32 r3263 (rst, clk, in, r3263_out);
	reg32 r3264 (rst, clk, in, r3264_out);
	reg32 r3265 (rst, clk, in, r3265_out);
	reg32 r3266 (rst, clk, in, r3266_out);
	reg32 r3267 (rst, clk, in, r3267_out);
	reg32 r3268 (rst, clk, in, r3268_out);
	reg32 r3269 (rst, clk, in, r3269_out);
	reg32 r3270 (rst, clk, in, r3270_out);
	reg32 r3271 (rst, clk, in, r3271_out);
	reg32 r3272 (rst, clk, in, r3272_out);
	reg32 r3273 (rst, clk, in, r3273_out);
	reg32 r3274 (rst, clk, in, r3274_out);
	reg32 r3275 (rst, clk, in, r3275_out);
	reg32 r3276 (rst, clk, in, r3276_out);
	reg32 r3277 (rst, clk, in, r3277_out);
	reg32 r3278 (rst, clk, in, r3278_out);
	reg32 r3279 (rst, clk, in, r3279_out);
	reg32 r3280 (rst, clk, in, r3280_out);
	reg32 r3281 (rst, clk, in, r3281_out);
	reg32 r3282 (rst, clk, in, r3282_out);
	reg32 r3283 (rst, clk, in, r3283_out);
	reg32 r3284 (rst, clk, in, r3284_out);
	reg32 r3285 (rst, clk, in, r3285_out);
	reg32 r3286 (rst, clk, in, r3286_out);
	reg32 r3287 (rst, clk, in, r3287_out);
	reg32 r3288 (rst, clk, in, r3288_out);
	reg32 r3289 (rst, clk, in, r3289_out);
	reg32 r3290 (rst, clk, in, r3290_out);
	reg32 r3291 (rst, clk, in, r3291_out);
	reg32 r3292 (rst, clk, in, r3292_out);
	reg32 r3293 (rst, clk, in, r3293_out);
	reg32 r3294 (rst, clk, in, r3294_out);
	reg32 r3295 (rst, clk, in, r3295_out);
	reg32 r3296 (rst, clk, in, r3296_out);
	reg32 r3297 (rst, clk, in, r3297_out);
	reg32 r3298 (rst, clk, in, r3298_out);
	reg32 r3299 (rst, clk, in, r3299_out);
	reg32 r3300 (rst, clk, in, r3300_out);
	reg32 r3301 (rst, clk, in, r3301_out);
	reg32 r3302 (rst, clk, in, r3302_out);
	reg32 r3303 (rst, clk, in, r3303_out);
	reg32 r3304 (rst, clk, in, r3304_out);
	reg32 r3305 (rst, clk, in, r3305_out);
	reg32 r3306 (rst, clk, in, r3306_out);
	reg32 r3307 (rst, clk, in, r3307_out);
	reg32 r3308 (rst, clk, in, r3308_out);
	reg32 r3309 (rst, clk, in, r3309_out);
	reg32 r3310 (rst, clk, in, r3310_out);
	reg32 r3311 (rst, clk, in, r3311_out);
	reg32 r3312 (rst, clk, in, r3312_out);
	reg32 r3313 (rst, clk, in, r3313_out);
	reg32 r3314 (rst, clk, in, r3314_out);
	reg32 r3315 (rst, clk, in, r3315_out);
	reg32 r3316 (rst, clk, in, r3316_out);
	reg32 r3317 (rst, clk, in, r3317_out);
	reg32 r3318 (rst, clk, in, r3318_out);
	reg32 r3319 (rst, clk, in, r3319_out);
	reg32 r3320 (rst, clk, in, r3320_out);
	reg32 r3321 (rst, clk, in, r3321_out);
	reg32 r3322 (rst, clk, in, r3322_out);
	reg32 r3323 (rst, clk, in, r3323_out);
	reg32 r3324 (rst, clk, in, r3324_out);
	reg32 r3325 (rst, clk, in, r3325_out);
	reg32 r3326 (rst, clk, in, r3326_out);
	reg32 r3327 (rst, clk, in, r3327_out);
	reg32 r3328 (rst, clk, in, r3328_out);
	reg32 r3329 (rst, clk, in, r3329_out);
	reg32 r3330 (rst, clk, in, r3330_out);
	reg32 r3331 (rst, clk, in, r3331_out);
	reg32 r3332 (rst, clk, in, r3332_out);
	reg32 r3333 (rst, clk, in, r3333_out);
	reg32 r3334 (rst, clk, in, r3334_out);
	reg32 r3335 (rst, clk, in, r3335_out);
	reg32 r3336 (rst, clk, in, r3336_out);
	reg32 r3337 (rst, clk, in, r3337_out);
	reg32 r3338 (rst, clk, in, r3338_out);
	reg32 r3339 (rst, clk, in, r3339_out);
	reg32 r3340 (rst, clk, in, r3340_out);
	reg32 r3341 (rst, clk, in, r3341_out);
	reg32 r3342 (rst, clk, in, r3342_out);
	reg32 r3343 (rst, clk, in, r3343_out);
	reg32 r3344 (rst, clk, in, r3344_out);
	reg32 r3345 (rst, clk, in, r3345_out);
	reg32 r3346 (rst, clk, in, r3346_out);
	reg32 r3347 (rst, clk, in, r3347_out);
	reg32 r3348 (rst, clk, in, r3348_out);
	reg32 r3349 (rst, clk, in, r3349_out);
	reg32 r3350 (rst, clk, in, r3350_out);
	reg32 r3351 (rst, clk, in, r3351_out);
	reg32 r3352 (rst, clk, in, r3352_out);
	reg32 r3353 (rst, clk, in, r3353_out);
	reg32 r3354 (rst, clk, in, r3354_out);
	reg32 r3355 (rst, clk, in, r3355_out);
	reg32 r3356 (rst, clk, in, r3356_out);
	reg32 r3357 (rst, clk, in, r3357_out);
	reg32 r3358 (rst, clk, in, r3358_out);
	reg32 r3359 (rst, clk, in, r3359_out);
	reg32 r3360 (rst, clk, in, r3360_out);
	reg32 r3361 (rst, clk, in, r3361_out);
	reg32 r3362 (rst, clk, in, r3362_out);
	reg32 r3363 (rst, clk, in, r3363_out);
	reg32 r3364 (rst, clk, in, r3364_out);
	reg32 r3365 (rst, clk, in, r3365_out);
	reg32 r3366 (rst, clk, in, r3366_out);
	reg32 r3367 (rst, clk, in, r3367_out);
	reg32 r3368 (rst, clk, in, r3368_out);
	reg32 r3369 (rst, clk, in, r3369_out);
	reg32 r3370 (rst, clk, in, r3370_out);
	reg32 r3371 (rst, clk, in, r3371_out);
	reg32 r3372 (rst, clk, in, r3372_out);
	reg32 r3373 (rst, clk, in, r3373_out);
	reg32 r3374 (rst, clk, in, r3374_out);
	reg32 r3375 (rst, clk, in, r3375_out);
	reg32 r3376 (rst, clk, in, r3376_out);
	reg32 r3377 (rst, clk, in, r3377_out);
	reg32 r3378 (rst, clk, in, r3378_out);
	reg32 r3379 (rst, clk, in, r3379_out);
	reg32 r3380 (rst, clk, in, r3380_out);
	reg32 r3381 (rst, clk, in, r3381_out);
	reg32 r3382 (rst, clk, in, r3382_out);
	reg32 r3383 (rst, clk, in, r3383_out);
	reg32 r3384 (rst, clk, in, r3384_out);
	reg32 r3385 (rst, clk, in, r3385_out);
	reg32 r3386 (rst, clk, in, r3386_out);
	reg32 r3387 (rst, clk, in, r3387_out);
	reg32 r3388 (rst, clk, in, r3388_out);
	reg32 r3389 (rst, clk, in, r3389_out);
	reg32 r3390 (rst, clk, in, r3390_out);
	reg32 r3391 (rst, clk, in, r3391_out);
	reg32 r3392 (rst, clk, in, r3392_out);
	reg32 r3393 (rst, clk, in, r3393_out);
	reg32 r3394 (rst, clk, in, r3394_out);
	reg32 r3395 (rst, clk, in, r3395_out);
	reg32 r3396 (rst, clk, in, r3396_out);
	reg32 r3397 (rst, clk, in, r3397_out);
	reg32 r3398 (rst, clk, in, r3398_out);
	reg32 r3399 (rst, clk, in, r3399_out);
	reg32 r3400 (rst, clk, in, r3400_out);
	reg32 r3401 (rst, clk, in, r3401_out);
	reg32 r3402 (rst, clk, in, r3402_out);
	reg32 r3403 (rst, clk, in, r3403_out);
	reg32 r3404 (rst, clk, in, r3404_out);
	reg32 r3405 (rst, clk, in, r3405_out);
	reg32 r3406 (rst, clk, in, r3406_out);
	reg32 r3407 (rst, clk, in, r3407_out);
	reg32 r3408 (rst, clk, in, r3408_out);
	reg32 r3409 (rst, clk, in, r3409_out);
	reg32 r3410 (rst, clk, in, r3410_out);
	reg32 r3411 (rst, clk, in, r3411_out);
	reg32 r3412 (rst, clk, in, r3412_out);
	reg32 r3413 (rst, clk, in, r3413_out);
	reg32 r3414 (rst, clk, in, r3414_out);
	reg32 r3415 (rst, clk, in, r3415_out);
	reg32 r3416 (rst, clk, in, r3416_out);
	reg32 r3417 (rst, clk, in, r3417_out);
	reg32 r3418 (rst, clk, in, r3418_out);
	reg32 r3419 (rst, clk, in, r3419_out);
	reg32 r3420 (rst, clk, in, r3420_out);
	reg32 r3421 (rst, clk, in, r3421_out);
	reg32 r3422 (rst, clk, in, r3422_out);
	reg32 r3423 (rst, clk, in, r3423_out);
	reg32 r3424 (rst, clk, in, r3424_out);
	reg32 r3425 (rst, clk, in, r3425_out);
	reg32 r3426 (rst, clk, in, r3426_out);
	reg32 r3427 (rst, clk, in, r3427_out);
	reg32 r3428 (rst, clk, in, r3428_out);
	reg32 r3429 (rst, clk, in, r3429_out);
	reg32 r3430 (rst, clk, in, r3430_out);
	reg32 r3431 (rst, clk, in, r3431_out);
	reg32 r3432 (rst, clk, in, r3432_out);
	reg32 r3433 (rst, clk, in, r3433_out);
	reg32 r3434 (rst, clk, in, r3434_out);
	reg32 r3435 (rst, clk, in, r3435_out);
	reg32 r3436 (rst, clk, in, r3436_out);
	reg32 r3437 (rst, clk, in, r3437_out);
	reg32 r3438 (rst, clk, in, r3438_out);
	reg32 r3439 (rst, clk, in, r3439_out);
	reg32 r3440 (rst, clk, in, r3440_out);
	reg32 r3441 (rst, clk, in, r3441_out);
	reg32 r3442 (rst, clk, in, r3442_out);
	reg32 r3443 (rst, clk, in, r3443_out);
	reg32 r3444 (rst, clk, in, r3444_out);
	reg32 r3445 (rst, clk, in, r3445_out);
	reg32 r3446 (rst, clk, in, r3446_out);
	reg32 r3447 (rst, clk, in, r3447_out);
	reg32 r3448 (rst, clk, in, r3448_out);
	reg32 r3449 (rst, clk, in, r3449_out);
	reg32 r3450 (rst, clk, in, r3450_out);
	reg32 r3451 (rst, clk, in, r3451_out);
	reg32 r3452 (rst, clk, in, r3452_out);
	reg32 r3453 (rst, clk, in, r3453_out);
	reg32 r3454 (rst, clk, in, r3454_out);
	reg32 r3455 (rst, clk, in, r3455_out);
	reg32 r3456 (rst, clk, in, r3456_out);
	reg32 r3457 (rst, clk, in, r3457_out);
	reg32 r3458 (rst, clk, in, r3458_out);
	reg32 r3459 (rst, clk, in, r3459_out);
	reg32 r3460 (rst, clk, in, r3460_out);
	reg32 r3461 (rst, clk, in, r3461_out);
	reg32 r3462 (rst, clk, in, r3462_out);
	reg32 r3463 (rst, clk, in, r3463_out);
	reg32 r3464 (rst, clk, in, r3464_out);
	reg32 r3465 (rst, clk, in, r3465_out);
	reg32 r3466 (rst, clk, in, r3466_out);
	reg32 r3467 (rst, clk, in, r3467_out);
	reg32 r3468 (rst, clk, in, r3468_out);
	reg32 r3469 (rst, clk, in, r3469_out);
	reg32 r3470 (rst, clk, in, r3470_out);
	reg32 r3471 (rst, clk, in, r3471_out);
	reg32 r3472 (rst, clk, in, r3472_out);
	reg32 r3473 (rst, clk, in, r3473_out);
	reg32 r3474 (rst, clk, in, r3474_out);
	reg32 r3475 (rst, clk, in, r3475_out);
	reg32 r3476 (rst, clk, in, r3476_out);
	reg32 r3477 (rst, clk, in, r3477_out);
	reg32 r3478 (rst, clk, in, r3478_out);
	reg32 r3479 (rst, clk, in, r3479_out);
	reg32 r3480 (rst, clk, in, r3480_out);
	reg32 r3481 (rst, clk, in, r3481_out);
	reg32 r3482 (rst, clk, in, r3482_out);
	reg32 r3483 (rst, clk, in, r3483_out);
	reg32 r3484 (rst, clk, in, r3484_out);
	reg32 r3485 (rst, clk, in, r3485_out);
	reg32 r3486 (rst, clk, in, r3486_out);
	reg32 r3487 (rst, clk, in, r3487_out);
	reg32 r3488 (rst, clk, in, r3488_out);
	reg32 r3489 (rst, clk, in, r3489_out);
	reg32 r3490 (rst, clk, in, r3490_out);
	reg32 r3491 (rst, clk, in, r3491_out);
	reg32 r3492 (rst, clk, in, r3492_out);
	reg32 r3493 (rst, clk, in, r3493_out);
	reg32 r3494 (rst, clk, in, r3494_out);
	reg32 r3495 (rst, clk, in, r3495_out);
	reg32 r3496 (rst, clk, in, r3496_out);
	reg32 r3497 (rst, clk, in, r3497_out);
	reg32 r3498 (rst, clk, in, r3498_out);
	reg32 r3499 (rst, clk, in, r3499_out);
	reg32 r3500 (rst, clk, in, r3500_out);
	reg32 r3501 (rst, clk, in, r3501_out);
	reg32 r3502 (rst, clk, in, r3502_out);
	reg32 r3503 (rst, clk, in, r3503_out);
	reg32 r3504 (rst, clk, in, r3504_out);
	reg32 r3505 (rst, clk, in, r3505_out);
	reg32 r3506 (rst, clk, in, r3506_out);
	reg32 r3507 (rst, clk, in, r3507_out);
	reg32 r3508 (rst, clk, in, r3508_out);
	reg32 r3509 (rst, clk, in, r3509_out);
	reg32 r3510 (rst, clk, in, r3510_out);
	reg32 r3511 (rst, clk, in, r3511_out);
	reg32 r3512 (rst, clk, in, r3512_out);
	reg32 r3513 (rst, clk, in, r3513_out);
	reg32 r3514 (rst, clk, in, r3514_out);
	reg32 r3515 (rst, clk, in, r3515_out);
	reg32 r3516 (rst, clk, in, r3516_out);
	reg32 r3517 (rst, clk, in, r3517_out);
	reg32 r3518 (rst, clk, in, r3518_out);
	reg32 r3519 (rst, clk, in, r3519_out);
	reg32 r3520 (rst, clk, in, r3520_out);
	reg32 r3521 (rst, clk, in, r3521_out);
	reg32 r3522 (rst, clk, in, r3522_out);
	reg32 r3523 (rst, clk, in, r3523_out);
	reg32 r3524 (rst, clk, in, r3524_out);
	reg32 r3525 (rst, clk, in, r3525_out);
	reg32 r3526 (rst, clk, in, r3526_out);
	reg32 r3527 (rst, clk, in, r3527_out);
	reg32 r3528 (rst, clk, in, r3528_out);
	reg32 r3529 (rst, clk, in, r3529_out);
	reg32 r3530 (rst, clk, in, r3530_out);
	reg32 r3531 (rst, clk, in, r3531_out);
	reg32 r3532 (rst, clk, in, r3532_out);
	reg32 r3533 (rst, clk, in, r3533_out);
	reg32 r3534 (rst, clk, in, r3534_out);
	reg32 r3535 (rst, clk, in, r3535_out);
	reg32 r3536 (rst, clk, in, r3536_out);
	reg32 r3537 (rst, clk, in, r3537_out);
	reg32 r3538 (rst, clk, in, r3538_out);
	reg32 r3539 (rst, clk, in, r3539_out);
	reg32 r3540 (rst, clk, in, r3540_out);
	reg32 r3541 (rst, clk, in, r3541_out);
	reg32 r3542 (rst, clk, in, r3542_out);
	reg32 r3543 (rst, clk, in, r3543_out);
	reg32 r3544 (rst, clk, in, r3544_out);
	reg32 r3545 (rst, clk, in, r3545_out);
	reg32 r3546 (rst, clk, in, r3546_out);
	reg32 r3547 (rst, clk, in, r3547_out);
	reg32 r3548 (rst, clk, in, r3548_out);
	reg32 r3549 (rst, clk, in, r3549_out);
	reg32 r3550 (rst, clk, in, r3550_out);
	reg32 r3551 (rst, clk, in, r3551_out);
	reg32 r3552 (rst, clk, in, r3552_out);
	reg32 r3553 (rst, clk, in, r3553_out);
	reg32 r3554 (rst, clk, in, r3554_out);
	reg32 r3555 (rst, clk, in, r3555_out);
	reg32 r3556 (rst, clk, in, r3556_out);
	reg32 r3557 (rst, clk, in, r3557_out);
	reg32 r3558 (rst, clk, in, r3558_out);
	reg32 r3559 (rst, clk, in, r3559_out);
	reg32 r3560 (rst, clk, in, r3560_out);
	reg32 r3561 (rst, clk, in, r3561_out);
	reg32 r3562 (rst, clk, in, r3562_out);
	reg32 r3563 (rst, clk, in, r3563_out);
	reg32 r3564 (rst, clk, in, r3564_out);
	reg32 r3565 (rst, clk, in, r3565_out);
	reg32 r3566 (rst, clk, in, r3566_out);
	reg32 r3567 (rst, clk, in, r3567_out);
	reg32 r3568 (rst, clk, in, r3568_out);
	reg32 r3569 (rst, clk, in, r3569_out);
	reg32 r3570 (rst, clk, in, r3570_out);
	reg32 r3571 (rst, clk, in, r3571_out);
	reg32 r3572 (rst, clk, in, r3572_out);
	reg32 r3573 (rst, clk, in, r3573_out);
	reg32 r3574 (rst, clk, in, r3574_out);
	reg32 r3575 (rst, clk, in, r3575_out);
	reg32 r3576 (rst, clk, in, r3576_out);
	reg32 r3577 (rst, clk, in, r3577_out);
	reg32 r3578 (rst, clk, in, r3578_out);
	reg32 r3579 (rst, clk, in, r3579_out);
	reg32 r3580 (rst, clk, in, r3580_out);
	reg32 r3581 (rst, clk, in, r3581_out);
	reg32 r3582 (rst, clk, in, r3582_out);
	reg32 r3583 (rst, clk, in, r3583_out);
	reg32 r3584 (rst, clk, in, r3584_out);
	reg32 r3585 (rst, clk, in, r3585_out);
	reg32 r3586 (rst, clk, in, r3586_out);
	reg32 r3587 (rst, clk, in, r3587_out);
	reg32 r3588 (rst, clk, in, r3588_out);
	reg32 r3589 (rst, clk, in, r3589_out);
	reg32 r3590 (rst, clk, in, r3590_out);
	reg32 r3591 (rst, clk, in, r3591_out);
	reg32 r3592 (rst, clk, in, r3592_out);
	reg32 r3593 (rst, clk, in, r3593_out);
	reg32 r3594 (rst, clk, in, r3594_out);
	reg32 r3595 (rst, clk, in, r3595_out);
	reg32 r3596 (rst, clk, in, r3596_out);
	reg32 r3597 (rst, clk, in, r3597_out);
	reg32 r3598 (rst, clk, in, r3598_out);
	reg32 r3599 (rst, clk, in, r3599_out);
	reg32 r3600 (rst, clk, in, r3600_out);
	reg32 r3601 (rst, clk, in, r3601_out);
	reg32 r3602 (rst, clk, in, r3602_out);
	reg32 r3603 (rst, clk, in, r3603_out);
	reg32 r3604 (rst, clk, in, r3604_out);
	reg32 r3605 (rst, clk, in, r3605_out);
	reg32 r3606 (rst, clk, in, r3606_out);
	reg32 r3607 (rst, clk, in, r3607_out);
	reg32 r3608 (rst, clk, in, r3608_out);
	reg32 r3609 (rst, clk, in, r3609_out);
	reg32 r3610 (rst, clk, in, r3610_out);
	reg32 r3611 (rst, clk, in, r3611_out);
	reg32 r3612 (rst, clk, in, r3612_out);
	reg32 r3613 (rst, clk, in, r3613_out);
	reg32 r3614 (rst, clk, in, r3614_out);
	reg32 r3615 (rst, clk, in, r3615_out);
	reg32 r3616 (rst, clk, in, r3616_out);
	reg32 r3617 (rst, clk, in, r3617_out);
	reg32 r3618 (rst, clk, in, r3618_out);
	reg32 r3619 (rst, clk, in, r3619_out);
	reg32 r3620 (rst, clk, in, r3620_out);
	reg32 r3621 (rst, clk, in, r3621_out);
	reg32 r3622 (rst, clk, in, r3622_out);
	reg32 r3623 (rst, clk, in, r3623_out);
	reg32 r3624 (rst, clk, in, r3624_out);
	reg32 r3625 (rst, clk, in, r3625_out);
	reg32 r3626 (rst, clk, in, r3626_out);
	reg32 r3627 (rst, clk, in, r3627_out);
	reg32 r3628 (rst, clk, in, r3628_out);
	reg32 r3629 (rst, clk, in, r3629_out);
	reg32 r3630 (rst, clk, in, r3630_out);
	reg32 r3631 (rst, clk, in, r3631_out);
	reg32 r3632 (rst, clk, in, r3632_out);
	reg32 r3633 (rst, clk, in, r3633_out);
	reg32 r3634 (rst, clk, in, r3634_out);
	reg32 r3635 (rst, clk, in, r3635_out);
	reg32 r3636 (rst, clk, in, r3636_out);
	reg32 r3637 (rst, clk, in, r3637_out);
	reg32 r3638 (rst, clk, in, r3638_out);
	reg32 r3639 (rst, clk, in, r3639_out);
	reg32 r3640 (rst, clk, in, r3640_out);
	reg32 r3641 (rst, clk, in, r3641_out);
	reg32 r3642 (rst, clk, in, r3642_out);
	reg32 r3643 (rst, clk, in, r3643_out);
	reg32 r3644 (rst, clk, in, r3644_out);
	reg32 r3645 (rst, clk, in, r3645_out);
	reg32 r3646 (rst, clk, in, r3646_out);
	reg32 r3647 (rst, clk, in, r3647_out);
	reg32 r3648 (rst, clk, in, r3648_out);
	reg32 r3649 (rst, clk, in, r3649_out);
	reg32 r3650 (rst, clk, in, r3650_out);
	reg32 r3651 (rst, clk, in, r3651_out);
	reg32 r3652 (rst, clk, in, r3652_out);
	reg32 r3653 (rst, clk, in, r3653_out);
	reg32 r3654 (rst, clk, in, r3654_out);
	reg32 r3655 (rst, clk, in, r3655_out);
	reg32 r3656 (rst, clk, in, r3656_out);
	reg32 r3657 (rst, clk, in, r3657_out);
	reg32 r3658 (rst, clk, in, r3658_out);
	reg32 r3659 (rst, clk, in, r3659_out);
	reg32 r3660 (rst, clk, in, r3660_out);
	reg32 r3661 (rst, clk, in, r3661_out);
	reg32 r3662 (rst, clk, in, r3662_out);
	reg32 r3663 (rst, clk, in, r3663_out);
	reg32 r3664 (rst, clk, in, r3664_out);
	reg32 r3665 (rst, clk, in, r3665_out);
	reg32 r3666 (rst, clk, in, r3666_out);
	reg32 r3667 (rst, clk, in, r3667_out);
	reg32 r3668 (rst, clk, in, r3668_out);
	reg32 r3669 (rst, clk, in, r3669_out);
	reg32 r3670 (rst, clk, in, r3670_out);
	reg32 r3671 (rst, clk, in, r3671_out);
	reg32 r3672 (rst, clk, in, r3672_out);
	reg32 r3673 (rst, clk, in, r3673_out);
	reg32 r3674 (rst, clk, in, r3674_out);
	reg32 r3675 (rst, clk, in, r3675_out);
	reg32 r3676 (rst, clk, in, r3676_out);
	reg32 r3677 (rst, clk, in, r3677_out);
	reg32 r3678 (rst, clk, in, r3678_out);
	reg32 r3679 (rst, clk, in, r3679_out);
	reg32 r3680 (rst, clk, in, r3680_out);
	reg32 r3681 (rst, clk, in, r3681_out);
	reg32 r3682 (rst, clk, in, r3682_out);
	reg32 r3683 (rst, clk, in, r3683_out);
	reg32 r3684 (rst, clk, in, r3684_out);
	reg32 r3685 (rst, clk, in, r3685_out);
	reg32 r3686 (rst, clk, in, r3686_out);
	reg32 r3687 (rst, clk, in, r3687_out);
	reg32 r3688 (rst, clk, in, r3688_out);
	reg32 r3689 (rst, clk, in, r3689_out);
	reg32 r3690 (rst, clk, in, r3690_out);
	reg32 r3691 (rst, clk, in, r3691_out);
	reg32 r3692 (rst, clk, in, r3692_out);
	reg32 r3693 (rst, clk, in, r3693_out);
	reg32 r3694 (rst, clk, in, r3694_out);
	reg32 r3695 (rst, clk, in, r3695_out);
	reg32 r3696 (rst, clk, in, r3696_out);
	reg32 r3697 (rst, clk, in, r3697_out);
	reg32 r3698 (rst, clk, in, r3698_out);
	reg32 r3699 (rst, clk, in, r3699_out);
	reg32 r3700 (rst, clk, in, r3700_out);
	reg32 r3701 (rst, clk, in, r3701_out);
	reg32 r3702 (rst, clk, in, r3702_out);
	reg32 r3703 (rst, clk, in, r3703_out);
	reg32 r3704 (rst, clk, in, r3704_out);
	reg32 r3705 (rst, clk, in, r3705_out);
	reg32 r3706 (rst, clk, in, r3706_out);
	reg32 r3707 (rst, clk, in, r3707_out);
	reg32 r3708 (rst, clk, in, r3708_out);
	reg32 r3709 (rst, clk, in, r3709_out);
	reg32 r3710 (rst, clk, in, r3710_out);
	reg32 r3711 (rst, clk, in, r3711_out);
	reg32 r3712 (rst, clk, in, r3712_out);
	reg32 r3713 (rst, clk, in, r3713_out);
	reg32 r3714 (rst, clk, in, r3714_out);
	reg32 r3715 (rst, clk, in, r3715_out);
	reg32 r3716 (rst, clk, in, r3716_out);
	reg32 r3717 (rst, clk, in, r3717_out);
	reg32 r3718 (rst, clk, in, r3718_out);
	reg32 r3719 (rst, clk, in, r3719_out);
	reg32 r3720 (rst, clk, in, r3720_out);
	reg32 r3721 (rst, clk, in, r3721_out);
	reg32 r3722 (rst, clk, in, r3722_out);
	reg32 r3723 (rst, clk, in, r3723_out);
	reg32 r3724 (rst, clk, in, r3724_out);
	reg32 r3725 (rst, clk, in, r3725_out);
	reg32 r3726 (rst, clk, in, r3726_out);
	reg32 r3727 (rst, clk, in, r3727_out);
	reg32 r3728 (rst, clk, in, r3728_out);
	reg32 r3729 (rst, clk, in, r3729_out);
	reg32 r3730 (rst, clk, in, r3730_out);
	reg32 r3731 (rst, clk, in, r3731_out);
	reg32 r3732 (rst, clk, in, r3732_out);
	reg32 r3733 (rst, clk, in, r3733_out);
	reg32 r3734 (rst, clk, in, r3734_out);
	reg32 r3735 (rst, clk, in, r3735_out);
	reg32 r3736 (rst, clk, in, r3736_out);
	reg32 r3737 (rst, clk, in, r3737_out);
	reg32 r3738 (rst, clk, in, r3738_out);
	reg32 r3739 (rst, clk, in, r3739_out);
	reg32 r3740 (rst, clk, in, r3740_out);
	reg32 r3741 (rst, clk, in, r3741_out);
	reg32 r3742 (rst, clk, in, r3742_out);
	reg32 r3743 (rst, clk, in, r3743_out);
	reg32 r3744 (rst, clk, in, r3744_out);
	reg32 r3745 (rst, clk, in, r3745_out);
	reg32 r3746 (rst, clk, in, r3746_out);
	reg32 r3747 (rst, clk, in, r3747_out);
	reg32 r3748 (rst, clk, in, r3748_out);
	reg32 r3749 (rst, clk, in, r3749_out);
	reg32 r3750 (rst, clk, in, r3750_out);
	reg32 r3751 (rst, clk, in, r3751_out);
	reg32 r3752 (rst, clk, in, r3752_out);
	reg32 r3753 (rst, clk, in, r3753_out);
	reg32 r3754 (rst, clk, in, r3754_out);
	reg32 r3755 (rst, clk, in, r3755_out);
	reg32 r3756 (rst, clk, in, r3756_out);
	reg32 r3757 (rst, clk, in, r3757_out);
	reg32 r3758 (rst, clk, in, r3758_out);
	reg32 r3759 (rst, clk, in, r3759_out);
	reg32 r3760 (rst, clk, in, r3760_out);
	reg32 r3761 (rst, clk, in, r3761_out);
	reg32 r3762 (rst, clk, in, r3762_out);
	reg32 r3763 (rst, clk, in, r3763_out);
	reg32 r3764 (rst, clk, in, r3764_out);
	reg32 r3765 (rst, clk, in, r3765_out);
	reg32 r3766 (rst, clk, in, r3766_out);
	reg32 r3767 (rst, clk, in, r3767_out);
	reg32 r3768 (rst, clk, in, r3768_out);
	reg32 r3769 (rst, clk, in, r3769_out);
	reg32 r3770 (rst, clk, in, r3770_out);
	reg32 r3771 (rst, clk, in, r3771_out);
	reg32 r3772 (rst, clk, in, r3772_out);
	reg32 r3773 (rst, clk, in, r3773_out);
	reg32 r3774 (rst, clk, in, r3774_out);
	reg32 r3775 (rst, clk, in, r3775_out);
	reg32 r3776 (rst, clk, in, r3776_out);
	reg32 r3777 (rst, clk, in, r3777_out);
	reg32 r3778 (rst, clk, in, r3778_out);
	reg32 r3779 (rst, clk, in, r3779_out);
	reg32 r3780 (rst, clk, in, r3780_out);
	reg32 r3781 (rst, clk, in, r3781_out);
	reg32 r3782 (rst, clk, in, r3782_out);
	reg32 r3783 (rst, clk, in, r3783_out);
	reg32 r3784 (rst, clk, in, r3784_out);
	reg32 r3785 (rst, clk, in, r3785_out);
	reg32 r3786 (rst, clk, in, r3786_out);
	reg32 r3787 (rst, clk, in, r3787_out);
	reg32 r3788 (rst, clk, in, r3788_out);
	reg32 r3789 (rst, clk, in, r3789_out);
	reg32 r3790 (rst, clk, in, r3790_out);
	reg32 r3791 (rst, clk, in, r3791_out);
	reg32 r3792 (rst, clk, in, r3792_out);
	reg32 r3793 (rst, clk, in, r3793_out);
	reg32 r3794 (rst, clk, in, r3794_out);
	reg32 r3795 (rst, clk, in, r3795_out);
	reg32 r3796 (rst, clk, in, r3796_out);
	reg32 r3797 (rst, clk, in, r3797_out);
	reg32 r3798 (rst, clk, in, r3798_out);
	reg32 r3799 (rst, clk, in, r3799_out);
	reg32 r3800 (rst, clk, in, r3800_out);
	reg32 r3801 (rst, clk, in, r3801_out);
	reg32 r3802 (rst, clk, in, r3802_out);
	reg32 r3803 (rst, clk, in, r3803_out);
	reg32 r3804 (rst, clk, in, r3804_out);
	reg32 r3805 (rst, clk, in, r3805_out);
	reg32 r3806 (rst, clk, in, r3806_out);
	reg32 r3807 (rst, clk, in, r3807_out);
	reg32 r3808 (rst, clk, in, r3808_out);
	reg32 r3809 (rst, clk, in, r3809_out);
	reg32 r3810 (rst, clk, in, r3810_out);
	reg32 r3811 (rst, clk, in, r3811_out);
	reg32 r3812 (rst, clk, in, r3812_out);
	reg32 r3813 (rst, clk, in, r3813_out);
	reg32 r3814 (rst, clk, in, r3814_out);
	reg32 r3815 (rst, clk, in, r3815_out);
	reg32 r3816 (rst, clk, in, r3816_out);
	reg32 r3817 (rst, clk, in, r3817_out);
	reg32 r3818 (rst, clk, in, r3818_out);
	reg32 r3819 (rst, clk, in, r3819_out);
	reg32 r3820 (rst, clk, in, r3820_out);
	reg32 r3821 (rst, clk, in, r3821_out);
	reg32 r3822 (rst, clk, in, r3822_out);
	reg32 r3823 (rst, clk, in, r3823_out);
	reg32 r3824 (rst, clk, in, r3824_out);
	reg32 r3825 (rst, clk, in, r3825_out);
	reg32 r3826 (rst, clk, in, r3826_out);
	reg32 r3827 (rst, clk, in, r3827_out);
	reg32 r3828 (rst, clk, in, r3828_out);
	reg32 r3829 (rst, clk, in, r3829_out);
	reg32 r3830 (rst, clk, in, r3830_out);
	reg32 r3831 (rst, clk, in, r3831_out);
	reg32 r3832 (rst, clk, in, r3832_out);
	reg32 r3833 (rst, clk, in, r3833_out);
	reg32 r3834 (rst, clk, in, r3834_out);
	reg32 r3835 (rst, clk, in, r3835_out);
	reg32 r3836 (rst, clk, in, r3836_out);
	reg32 r3837 (rst, clk, in, r3837_out);
	reg32 r3838 (rst, clk, in, r3838_out);
	reg32 r3839 (rst, clk, in, r3839_out);
	reg32 r3840 (rst, clk, in, r3840_out);
	reg32 r3841 (rst, clk, in, r3841_out);
	reg32 r3842 (rst, clk, in, r3842_out);
	reg32 r3843 (rst, clk, in, r3843_out);
	reg32 r3844 (rst, clk, in, r3844_out);
	reg32 r3845 (rst, clk, in, r3845_out);
	reg32 r3846 (rst, clk, in, r3846_out);
	reg32 r3847 (rst, clk, in, r3847_out);
	reg32 r3848 (rst, clk, in, r3848_out);
	reg32 r3849 (rst, clk, in, r3849_out);
	reg32 r3850 (rst, clk, in, r3850_out);
	reg32 r3851 (rst, clk, in, r3851_out);
	reg32 r3852 (rst, clk, in, r3852_out);
	reg32 r3853 (rst, clk, in, r3853_out);
	reg32 r3854 (rst, clk, in, r3854_out);
	reg32 r3855 (rst, clk, in, r3855_out);
	reg32 r3856 (rst, clk, in, r3856_out);
	reg32 r3857 (rst, clk, in, r3857_out);
	reg32 r3858 (rst, clk, in, r3858_out);
	reg32 r3859 (rst, clk, in, r3859_out);
	reg32 r3860 (rst, clk, in, r3860_out);
	reg32 r3861 (rst, clk, in, r3861_out);
	reg32 r3862 (rst, clk, in, r3862_out);
	reg32 r3863 (rst, clk, in, r3863_out);
	reg32 r3864 (rst, clk, in, r3864_out);
	reg32 r3865 (rst, clk, in, r3865_out);
	reg32 r3866 (rst, clk, in, r3866_out);
	reg32 r3867 (rst, clk, in, r3867_out);
	reg32 r3868 (rst, clk, in, r3868_out);
	reg32 r3869 (rst, clk, in, r3869_out);
	reg32 r3870 (rst, clk, in, r3870_out);
	reg32 r3871 (rst, clk, in, r3871_out);
	reg32 r3872 (rst, clk, in, r3872_out);
	reg32 r3873 (rst, clk, in, r3873_out);
	reg32 r3874 (rst, clk, in, r3874_out);
	reg32 r3875 (rst, clk, in, r3875_out);
	reg32 r3876 (rst, clk, in, r3876_out);
	reg32 r3877 (rst, clk, in, r3877_out);
	reg32 r3878 (rst, clk, in, r3878_out);
	reg32 r3879 (rst, clk, in, r3879_out);
	reg32 r3880 (rst, clk, in, r3880_out);
	reg32 r3881 (rst, clk, in, r3881_out);
	reg32 r3882 (rst, clk, in, r3882_out);
	reg32 r3883 (rst, clk, in, r3883_out);
	reg32 r3884 (rst, clk, in, r3884_out);
	reg32 r3885 (rst, clk, in, r3885_out);
	reg32 r3886 (rst, clk, in, r3886_out);
	reg32 r3887 (rst, clk, in, r3887_out);
	reg32 r3888 (rst, clk, in, r3888_out);
	reg32 r3889 (rst, clk, in, r3889_out);
	reg32 r3890 (rst, clk, in, r3890_out);
	reg32 r3891 (rst, clk, in, r3891_out);
	reg32 r3892 (rst, clk, in, r3892_out);
	reg32 r3893 (rst, clk, in, r3893_out);
	reg32 r3894 (rst, clk, in, r3894_out);
	reg32 r3895 (rst, clk, in, r3895_out);
	reg32 r3896 (rst, clk, in, r3896_out);
	reg32 r3897 (rst, clk, in, r3897_out);
	reg32 r3898 (rst, clk, in, r3898_out);
	reg32 r3899 (rst, clk, in, r3899_out);
	reg32 r3900 (rst, clk, in, r3900_out);
	reg32 r3901 (rst, clk, in, r3901_out);
	reg32 r3902 (rst, clk, in, r3902_out);
	reg32 r3903 (rst, clk, in, r3903_out);
	reg32 r3904 (rst, clk, in, r3904_out);
	reg32 r3905 (rst, clk, in, r3905_out);
	reg32 r3906 (rst, clk, in, r3906_out);
	reg32 r3907 (rst, clk, in, r3907_out);
	reg32 r3908 (rst, clk, in, r3908_out);
	reg32 r3909 (rst, clk, in, r3909_out);
	reg32 r3910 (rst, clk, in, r3910_out);
	reg32 r3911 (rst, clk, in, r3911_out);
	reg32 r3912 (rst, clk, in, r3912_out);
	reg32 r3913 (rst, clk, in, r3913_out);
	reg32 r3914 (rst, clk, in, r3914_out);
	reg32 r3915 (rst, clk, in, r3915_out);
	reg32 r3916 (rst, clk, in, r3916_out);
	reg32 r3917 (rst, clk, in, r3917_out);
	reg32 r3918 (rst, clk, in, r3918_out);
	reg32 r3919 (rst, clk, in, r3919_out);
	reg32 r3920 (rst, clk, in, r3920_out);
	reg32 r3921 (rst, clk, in, r3921_out);
	reg32 r3922 (rst, clk, in, r3922_out);
	reg32 r3923 (rst, clk, in, r3923_out);
	reg32 r3924 (rst, clk, in, r3924_out);
	reg32 r3925 (rst, clk, in, r3925_out);
	reg32 r3926 (rst, clk, in, r3926_out);
	reg32 r3927 (rst, clk, in, r3927_out);
	reg32 r3928 (rst, clk, in, r3928_out);
	reg32 r3929 (rst, clk, in, r3929_out);
	reg32 r3930 (rst, clk, in, r3930_out);
	reg32 r3931 (rst, clk, in, r3931_out);
	reg32 r3932 (rst, clk, in, r3932_out);
	reg32 r3933 (rst, clk, in, r3933_out);
	reg32 r3934 (rst, clk, in, r3934_out);
	reg32 r3935 (rst, clk, in, r3935_out);
	reg32 r3936 (rst, clk, in, r3936_out);
	reg32 r3937 (rst, clk, in, r3937_out);
	reg32 r3938 (rst, clk, in, r3938_out);
	reg32 r3939 (rst, clk, in, r3939_out);
	reg32 r3940 (rst, clk, in, r3940_out);
	reg32 r3941 (rst, clk, in, r3941_out);
	reg32 r3942 (rst, clk, in, r3942_out);
	reg32 r3943 (rst, clk, in, r3943_out);
	reg32 r3944 (rst, clk, in, r3944_out);
	reg32 r3945 (rst, clk, in, r3945_out);
	reg32 r3946 (rst, clk, in, r3946_out);
	reg32 r3947 (rst, clk, in, r3947_out);
	reg32 r3948 (rst, clk, in, r3948_out);
	reg32 r3949 (rst, clk, in, r3949_out);
	reg32 r3950 (rst, clk, in, r3950_out);
	reg32 r3951 (rst, clk, in, r3951_out);
	reg32 r3952 (rst, clk, in, r3952_out);
	reg32 r3953 (rst, clk, in, r3953_out);
	reg32 r3954 (rst, clk, in, r3954_out);
	reg32 r3955 (rst, clk, in, r3955_out);
	reg32 r3956 (rst, clk, in, r3956_out);
	reg32 r3957 (rst, clk, in, r3957_out);
	reg32 r3958 (rst, clk, in, r3958_out);
	reg32 r3959 (rst, clk, in, r3959_out);
	reg32 r3960 (rst, clk, in, r3960_out);
	reg32 r3961 (rst, clk, in, r3961_out);
	reg32 r3962 (rst, clk, in, r3962_out);
	reg32 r3963 (rst, clk, in, r3963_out);
	reg32 r3964 (rst, clk, in, r3964_out);
	reg32 r3965 (rst, clk, in, r3965_out);
	reg32 r3966 (rst, clk, in, r3966_out);
	reg32 r3967 (rst, clk, in, r3967_out);
	reg32 r3968 (rst, clk, in, r3968_out);
	reg32 r3969 (rst, clk, in, r3969_out);
	reg32 r3970 (rst, clk, in, r3970_out);
	reg32 r3971 (rst, clk, in, r3971_out);
	reg32 r3972 (rst, clk, in, r3972_out);
	reg32 r3973 (rst, clk, in, r3973_out);
	reg32 r3974 (rst, clk, in, r3974_out);
	reg32 r3975 (rst, clk, in, r3975_out);
	reg32 r3976 (rst, clk, in, r3976_out);
	reg32 r3977 (rst, clk, in, r3977_out);
	reg32 r3978 (rst, clk, in, r3978_out);
	reg32 r3979 (rst, clk, in, r3979_out);
	reg32 r3980 (rst, clk, in, r3980_out);
	reg32 r3981 (rst, clk, in, r3981_out);
	reg32 r3982 (rst, clk, in, r3982_out);
	reg32 r3983 (rst, clk, in, r3983_out);
	reg32 r3984 (rst, clk, in, r3984_out);
	reg32 r3985 (rst, clk, in, r3985_out);
	reg32 r3986 (rst, clk, in, r3986_out);
	reg32 r3987 (rst, clk, in, r3987_out);
	reg32 r3988 (rst, clk, in, r3988_out);
	reg32 r3989 (rst, clk, in, r3989_out);
	reg32 r3990 (rst, clk, in, r3990_out);
	reg32 r3991 (rst, clk, in, r3991_out);
	reg32 r3992 (rst, clk, in, r3992_out);
	reg32 r3993 (rst, clk, in, r3993_out);
	reg32 r3994 (rst, clk, in, r3994_out);
	reg32 r3995 (rst, clk, in, r3995_out);
	reg32 r3996 (rst, clk, in, r3996_out);
	reg32 r3997 (rst, clk, in, r3997_out);
	reg32 r3998 (rst, clk, in, r3998_out);
	reg32 r3999 (rst, clk, in, r3999_out);
	reg32 r4000 (rst, clk, in, r4000_out);
	reg32 r4001 (rst, clk, in, r4001_out);
	reg32 r4002 (rst, clk, in, r4002_out);
	reg32 r4003 (rst, clk, in, r4003_out);
	reg32 r4004 (rst, clk, in, r4004_out);
	reg32 r4005 (rst, clk, in, r4005_out);
	reg32 r4006 (rst, clk, in, r4006_out);
	reg32 r4007 (rst, clk, in, r4007_out);
	reg32 r4008 (rst, clk, in, r4008_out);
	reg32 r4009 (rst, clk, in, r4009_out);
	reg32 r4010 (rst, clk, in, r4010_out);
	reg32 r4011 (rst, clk, in, r4011_out);
	reg32 r4012 (rst, clk, in, r4012_out);
	reg32 r4013 (rst, clk, in, r4013_out);
	reg32 r4014 (rst, clk, in, r4014_out);
	reg32 r4015 (rst, clk, in, r4015_out);
	reg32 r4016 (rst, clk, in, r4016_out);
	reg32 r4017 (rst, clk, in, r4017_out);
	reg32 r4018 (rst, clk, in, r4018_out);
	reg32 r4019 (rst, clk, in, r4019_out);
	reg32 r4020 (rst, clk, in, r4020_out);
	reg32 r4021 (rst, clk, in, r4021_out);
	reg32 r4022 (rst, clk, in, r4022_out);
	reg32 r4023 (rst, clk, in, r4023_out);
	reg32 r4024 (rst, clk, in, r4024_out);
	reg32 r4025 (rst, clk, in, r4025_out);
	reg32 r4026 (rst, clk, in, r4026_out);
	reg32 r4027 (rst, clk, in, r4027_out);
	reg32 r4028 (rst, clk, in, r4028_out);
	reg32 r4029 (rst, clk, in, r4029_out);
	reg32 r4030 (rst, clk, in, r4030_out);
	reg32 r4031 (rst, clk, in, r4031_out);
	reg32 r4032 (rst, clk, in, r4032_out);
	reg32 r4033 (rst, clk, in, r4033_out);
	reg32 r4034 (rst, clk, in, r4034_out);
	reg32 r4035 (rst, clk, in, r4035_out);
	reg32 r4036 (rst, clk, in, r4036_out);
	reg32 r4037 (rst, clk, in, r4037_out);
	reg32 r4038 (rst, clk, in, r4038_out);
	reg32 r4039 (rst, clk, in, r4039_out);
	reg32 r4040 (rst, clk, in, r4040_out);
	reg32 r4041 (rst, clk, in, r4041_out);
	reg32 r4042 (rst, clk, in, r4042_out);
	reg32 r4043 (rst, clk, in, r4043_out);
	reg32 r4044 (rst, clk, in, r4044_out);
	reg32 r4045 (rst, clk, in, r4045_out);
	reg32 r4046 (rst, clk, in, r4046_out);
	reg32 r4047 (rst, clk, in, r4047_out);
	reg32 r4048 (rst, clk, in, r4048_out);
	reg32 r4049 (rst, clk, in, r4049_out);
	reg32 r4050 (rst, clk, in, r4050_out);
	reg32 r4051 (rst, clk, in, r4051_out);
	reg32 r4052 (rst, clk, in, r4052_out);
	reg32 r4053 (rst, clk, in, r4053_out);
	reg32 r4054 (rst, clk, in, r4054_out);
	reg32 r4055 (rst, clk, in, r4055_out);
	reg32 r4056 (rst, clk, in, r4056_out);
	reg32 r4057 (rst, clk, in, r4057_out);
	reg32 r4058 (rst, clk, in, r4058_out);
	reg32 r4059 (rst, clk, in, r4059_out);
	reg32 r4060 (rst, clk, in, r4060_out);
	reg32 r4061 (rst, clk, in, r4061_out);
	reg32 r4062 (rst, clk, in, r4062_out);
	reg32 r4063 (rst, clk, in, r4063_out);
	reg32 r4064 (rst, clk, in, r4064_out);
	reg32 r4065 (rst, clk, in, r4065_out);
	reg32 r4066 (rst, clk, in, r4066_out);
	reg32 r4067 (rst, clk, in, r4067_out);
	reg32 r4068 (rst, clk, in, r4068_out);
	reg32 r4069 (rst, clk, in, r4069_out);
	reg32 r4070 (rst, clk, in, r4070_out);
	reg32 r4071 (rst, clk, in, r4071_out);
	reg32 r4072 (rst, clk, in, r4072_out);
	reg32 r4073 (rst, clk, in, r4073_out);
	reg32 r4074 (rst, clk, in, r4074_out);
	reg32 r4075 (rst, clk, in, r4075_out);
	reg32 r4076 (rst, clk, in, r4076_out);
	reg32 r4077 (rst, clk, in, r4077_out);
	reg32 r4078 (rst, clk, in, r4078_out);
	reg32 r4079 (rst, clk, in, r4079_out);
	reg32 r4080 (rst, clk, in, r4080_out);
	reg32 r4081 (rst, clk, in, r4081_out);
	reg32 r4082 (rst, clk, in, r4082_out);
	reg32 r4083 (rst, clk, in, r4083_out);
	reg32 r4084 (rst, clk, in, r4084_out);
	reg32 r4085 (rst, clk, in, r4085_out);
	reg32 r4086 (rst, clk, in, r4086_out);
	reg32 r4087 (rst, clk, in, r4087_out);
	reg32 r4088 (rst, clk, in, r4088_out);
	reg32 r4089 (rst, clk, in, r4089_out);
	reg32 r4090 (rst, clk, in, r4090_out);
	reg32 r4091 (rst, clk, in, r4091_out);
	reg32 r4092 (rst, clk, in, r4092_out);
	reg32 r4093 (rst, clk, in, r4093_out);
	reg32 r4094 (rst, clk, in, r4094_out);
	reg32 r4095 (rst, clk, in, r4095_out);
	reg32 r4096 (rst, clk, in, r4096_out);
	reg32 r4097 (rst, clk, in, r4097_out);
	reg32 r4098 (rst, clk, in, r4098_out);
	reg32 r4099 (rst, clk, in, r4099_out);
	reg32 r4100 (rst, clk, in, r4100_out);
	reg32 r4101 (rst, clk, in, r4101_out);
	reg32 r4102 (rst, clk, in, r4102_out);
	reg32 r4103 (rst, clk, in, r4103_out);
	reg32 r4104 (rst, clk, in, r4104_out);
	reg32 r4105 (rst, clk, in, r4105_out);
	reg32 r4106 (rst, clk, in, r4106_out);
	reg32 r4107 (rst, clk, in, r4107_out);
	reg32 r4108 (rst, clk, in, r4108_out);
	reg32 r4109 (rst, clk, in, r4109_out);
	reg32 r4110 (rst, clk, in, r4110_out);
	reg32 r4111 (rst, clk, in, r4111_out);
	reg32 r4112 (rst, clk, in, r4112_out);
	reg32 r4113 (rst, clk, in, r4113_out);
	reg32 r4114 (rst, clk, in, r4114_out);
	reg32 r4115 (rst, clk, in, r4115_out);
	reg32 r4116 (rst, clk, in, r4116_out);
	reg32 r4117 (rst, clk, in, r4117_out);
	reg32 r4118 (rst, clk, in, r4118_out);
	reg32 r4119 (rst, clk, in, r4119_out);
	reg32 r4120 (rst, clk, in, r4120_out);
	reg32 r4121 (rst, clk, in, r4121_out);
	reg32 r4122 (rst, clk, in, r4122_out);
	reg32 r4123 (rst, clk, in, r4123_out);
	reg32 r4124 (rst, clk, in, r4124_out);
	reg32 r4125 (rst, clk, in, r4125_out);
	reg32 r4126 (rst, clk, in, r4126_out);
	reg32 r4127 (rst, clk, in, r4127_out);
	reg32 r4128 (rst, clk, in, r4128_out);
	reg32 r4129 (rst, clk, in, r4129_out);
	reg32 r4130 (rst, clk, in, r4130_out);
	reg32 r4131 (rst, clk, in, r4131_out);
	reg32 r4132 (rst, clk, in, r4132_out);
	reg32 r4133 (rst, clk, in, r4133_out);
	reg32 r4134 (rst, clk, in, r4134_out);
	reg32 r4135 (rst, clk, in, r4135_out);
	reg32 r4136 (rst, clk, in, r4136_out);
	reg32 r4137 (rst, clk, in, r4137_out);
	reg32 r4138 (rst, clk, in, r4138_out);
	reg32 r4139 (rst, clk, in, r4139_out);
	reg32 r4140 (rst, clk, in, r4140_out);
	reg32 r4141 (rst, clk, in, r4141_out);
	reg32 r4142 (rst, clk, in, r4142_out);
	reg32 r4143 (rst, clk, in, r4143_out);
	reg32 r4144 (rst, clk, in, r4144_out);
	reg32 r4145 (rst, clk, in, r4145_out);
	reg32 r4146 (rst, clk, in, r4146_out);
	reg32 r4147 (rst, clk, in, r4147_out);
	reg32 r4148 (rst, clk, in, r4148_out);
	reg32 r4149 (rst, clk, in, r4149_out);
	reg32 r4150 (rst, clk, in, r4150_out);
	reg32 r4151 (rst, clk, in, r4151_out);
	reg32 r4152 (rst, clk, in, r4152_out);
	reg32 r4153 (rst, clk, in, r4153_out);
	reg32 r4154 (rst, clk, in, r4154_out);
	reg32 r4155 (rst, clk, in, r4155_out);
	reg32 r4156 (rst, clk, in, r4156_out);
	reg32 r4157 (rst, clk, in, r4157_out);
	reg32 r4158 (rst, clk, in, r4158_out);
	reg32 r4159 (rst, clk, in, r4159_out);
	reg32 r4160 (rst, clk, in, r4160_out);
	reg32 r4161 (rst, clk, in, r4161_out);
	reg32 r4162 (rst, clk, in, r4162_out);
	reg32 r4163 (rst, clk, in, r4163_out);
	reg32 r4164 (rst, clk, in, r4164_out);
	reg32 r4165 (rst, clk, in, r4165_out);
	reg32 r4166 (rst, clk, in, r4166_out);
	reg32 r4167 (rst, clk, in, r4167_out);
	reg32 r4168 (rst, clk, in, r4168_out);
	reg32 r4169 (rst, clk, in, r4169_out);
	reg32 r4170 (rst, clk, in, r4170_out);
	reg32 r4171 (rst, clk, in, r4171_out);
	reg32 r4172 (rst, clk, in, r4172_out);
	reg32 r4173 (rst, clk, in, r4173_out);
	reg32 r4174 (rst, clk, in, r4174_out);
	reg32 r4175 (rst, clk, in, r4175_out);
	reg32 r4176 (rst, clk, in, r4176_out);
	reg32 r4177 (rst, clk, in, r4177_out);
	reg32 r4178 (rst, clk, in, r4178_out);
	reg32 r4179 (rst, clk, in, r4179_out);
	reg32 r4180 (rst, clk, in, r4180_out);
	reg32 r4181 (rst, clk, in, r4181_out);
	reg32 r4182 (rst, clk, in, r4182_out);
	reg32 r4183 (rst, clk, in, r4183_out);
	reg32 r4184 (rst, clk, in, r4184_out);
	reg32 r4185 (rst, clk, in, r4185_out);
	reg32 r4186 (rst, clk, in, r4186_out);
	reg32 r4187 (rst, clk, in, r4187_out);
	reg32 r4188 (rst, clk, in, r4188_out);
	reg32 r4189 (rst, clk, in, r4189_out);
	reg32 r4190 (rst, clk, in, r4190_out);
	reg32 r4191 (rst, clk, in, r4191_out);
	reg32 r4192 (rst, clk, in, r4192_out);
	reg32 r4193 (rst, clk, in, r4193_out);
	reg32 r4194 (rst, clk, in, r4194_out);
	reg32 r4195 (rst, clk, in, r4195_out);
	reg32 r4196 (rst, clk, in, r4196_out);
	reg32 r4197 (rst, clk, in, r4197_out);
	reg32 r4198 (rst, clk, in, r4198_out);
	reg32 r4199 (rst, clk, in, r4199_out);
	reg32 r4200 (rst, clk, in, r4200_out);
	reg32 r4201 (rst, clk, in, r4201_out);
	reg32 r4202 (rst, clk, in, r4202_out);
	reg32 r4203 (rst, clk, in, r4203_out);
	reg32 r4204 (rst, clk, in, r4204_out);
	reg32 r4205 (rst, clk, in, r4205_out);
	reg32 r4206 (rst, clk, in, r4206_out);
	reg32 r4207 (rst, clk, in, r4207_out);
	reg32 r4208 (rst, clk, in, r4208_out);
	reg32 r4209 (rst, clk, in, r4209_out);
	reg32 r4210 (rst, clk, in, r4210_out);
	reg32 r4211 (rst, clk, in, r4211_out);
	reg32 r4212 (rst, clk, in, r4212_out);
	reg32 r4213 (rst, clk, in, r4213_out);
	reg32 r4214 (rst, clk, in, r4214_out);
	reg32 r4215 (rst, clk, in, r4215_out);
	reg32 r4216 (rst, clk, in, r4216_out);
	reg32 r4217 (rst, clk, in, r4217_out);
	reg32 r4218 (rst, clk, in, r4218_out);
	reg32 r4219 (rst, clk, in, r4219_out);
	reg32 r4220 (rst, clk, in, r4220_out);
	reg32 r4221 (rst, clk, in, r4221_out);
	reg32 r4222 (rst, clk, in, r4222_out);
	reg32 r4223 (rst, clk, in, r4223_out);
	reg32 r4224 (rst, clk, in, r4224_out);
	reg32 r4225 (rst, clk, in, r4225_out);
	reg32 r4226 (rst, clk, in, r4226_out);
	reg32 r4227 (rst, clk, in, r4227_out);
	reg32 r4228 (rst, clk, in, r4228_out);
	reg32 r4229 (rst, clk, in, r4229_out);
	reg32 r4230 (rst, clk, in, r4230_out);
	reg32 r4231 (rst, clk, in, r4231_out);
	reg32 r4232 (rst, clk, in, r4232_out);
	reg32 r4233 (rst, clk, in, r4233_out);
	reg32 r4234 (rst, clk, in, r4234_out);
	reg32 r4235 (rst, clk, in, r4235_out);
	reg32 r4236 (rst, clk, in, r4236_out);
	reg32 r4237 (rst, clk, in, r4237_out);
	reg32 r4238 (rst, clk, in, r4238_out);
	reg32 r4239 (rst, clk, in, r4239_out);
	reg32 r4240 (rst, clk, in, r4240_out);
	reg32 r4241 (rst, clk, in, r4241_out);
	reg32 r4242 (rst, clk, in, r4242_out);
	reg32 r4243 (rst, clk, in, r4243_out);
	reg32 r4244 (rst, clk, in, r4244_out);
	reg32 r4245 (rst, clk, in, r4245_out);
	reg32 r4246 (rst, clk, in, r4246_out);
	reg32 r4247 (rst, clk, in, r4247_out);
	reg32 r4248 (rst, clk, in, r4248_out);
	reg32 r4249 (rst, clk, in, r4249_out);
	reg32 r4250 (rst, clk, in, r4250_out);
	reg32 r4251 (rst, clk, in, r4251_out);
	reg32 r4252 (rst, clk, in, r4252_out);
	reg32 r4253 (rst, clk, in, r4253_out);
	reg32 r4254 (rst, clk, in, r4254_out);
	reg32 r4255 (rst, clk, in, r4255_out);
	reg32 r4256 (rst, clk, in, r4256_out);
	reg32 r4257 (rst, clk, in, r4257_out);
	reg32 r4258 (rst, clk, in, r4258_out);
	reg32 r4259 (rst, clk, in, r4259_out);
	reg32 r4260 (rst, clk, in, r4260_out);
	reg32 r4261 (rst, clk, in, r4261_out);
	reg32 r4262 (rst, clk, in, r4262_out);
	reg32 r4263 (rst, clk, in, r4263_out);
	reg32 r4264 (rst, clk, in, r4264_out);
	reg32 r4265 (rst, clk, in, r4265_out);
	reg32 r4266 (rst, clk, in, r4266_out);
	reg32 r4267 (rst, clk, in, r4267_out);
	reg32 r4268 (rst, clk, in, r4268_out);
	reg32 r4269 (rst, clk, in, r4269_out);
	reg32 r4270 (rst, clk, in, r4270_out);
	reg32 r4271 (rst, clk, in, r4271_out);
	reg32 r4272 (rst, clk, in, r4272_out);
	reg32 r4273 (rst, clk, in, r4273_out);
	reg32 r4274 (rst, clk, in, r4274_out);
	reg32 r4275 (rst, clk, in, r4275_out);
	reg32 r4276 (rst, clk, in, r4276_out);
	reg32 r4277 (rst, clk, in, r4277_out);
	reg32 r4278 (rst, clk, in, r4278_out);
	reg32 r4279 (rst, clk, in, r4279_out);
	reg32 r4280 (rst, clk, in, r4280_out);
	reg32 r4281 (rst, clk, in, r4281_out);
	reg32 r4282 (rst, clk, in, r4282_out);
	reg32 r4283 (rst, clk, in, r4283_out);
	reg32 r4284 (rst, clk, in, r4284_out);
	reg32 r4285 (rst, clk, in, r4285_out);
	reg32 r4286 (rst, clk, in, r4286_out);
	reg32 r4287 (rst, clk, in, r4287_out);
	reg32 r4288 (rst, clk, in, r4288_out);
	reg32 r4289 (rst, clk, in, r4289_out);
	reg32 r4290 (rst, clk, in, r4290_out);
	reg32 r4291 (rst, clk, in, r4291_out);
	reg32 r4292 (rst, clk, in, r4292_out);
	reg32 r4293 (rst, clk, in, r4293_out);
	reg32 r4294 (rst, clk, in, r4294_out);
	reg32 r4295 (rst, clk, in, r4295_out);
	reg32 r4296 (rst, clk, in, r4296_out);
	reg32 r4297 (rst, clk, in, r4297_out);
	reg32 r4298 (rst, clk, in, r4298_out);
	reg32 r4299 (rst, clk, in, r4299_out);
	reg32 r4300 (rst, clk, in, r4300_out);
	reg32 r4301 (rst, clk, in, r4301_out);
	reg32 r4302 (rst, clk, in, r4302_out);
	reg32 r4303 (rst, clk, in, r4303_out);
	reg32 r4304 (rst, clk, in, r4304_out);
	reg32 r4305 (rst, clk, in, r4305_out);
	reg32 r4306 (rst, clk, in, r4306_out);
	reg32 r4307 (rst, clk, in, r4307_out);
	reg32 r4308 (rst, clk, in, r4308_out);
	reg32 r4309 (rst, clk, in, r4309_out);
	reg32 r4310 (rst, clk, in, r4310_out);
	reg32 r4311 (rst, clk, in, r4311_out);
	reg32 r4312 (rst, clk, in, r4312_out);
	reg32 r4313 (rst, clk, in, r4313_out);
	reg32 r4314 (rst, clk, in, r4314_out);
	reg32 r4315 (rst, clk, in, r4315_out);
	reg32 r4316 (rst, clk, in, r4316_out);
	reg32 r4317 (rst, clk, in, r4317_out);
	reg32 r4318 (rst, clk, in, r4318_out);
	reg32 r4319 (rst, clk, in, r4319_out);
	reg32 r4320 (rst, clk, in, r4320_out);
	reg32 r4321 (rst, clk, in, r4321_out);
	reg32 r4322 (rst, clk, in, r4322_out);
	reg32 r4323 (rst, clk, in, r4323_out);
	reg32 r4324 (rst, clk, in, r4324_out);
	reg32 r4325 (rst, clk, in, r4325_out);
	reg32 r4326 (rst, clk, in, r4326_out);
	reg32 r4327 (rst, clk, in, r4327_out);
	reg32 r4328 (rst, clk, in, r4328_out);
	reg32 r4329 (rst, clk, in, r4329_out);
	reg32 r4330 (rst, clk, in, r4330_out);
	reg32 r4331 (rst, clk, in, r4331_out);
	reg32 r4332 (rst, clk, in, r4332_out);
	reg32 r4333 (rst, clk, in, r4333_out);
	reg32 r4334 (rst, clk, in, r4334_out);
	reg32 r4335 (rst, clk, in, r4335_out);
	reg32 r4336 (rst, clk, in, r4336_out);
	reg32 r4337 (rst, clk, in, r4337_out);
	reg32 r4338 (rst, clk, in, r4338_out);
	reg32 r4339 (rst, clk, in, r4339_out);
	reg32 r4340 (rst, clk, in, r4340_out);
	reg32 r4341 (rst, clk, in, r4341_out);
	reg32 r4342 (rst, clk, in, r4342_out);
	reg32 r4343 (rst, clk, in, r4343_out);
	reg32 r4344 (rst, clk, in, r4344_out);
	reg32 r4345 (rst, clk, in, r4345_out);
	reg32 r4346 (rst, clk, in, r4346_out);
	reg32 r4347 (rst, clk, in, r4347_out);
	reg32 r4348 (rst, clk, in, r4348_out);
	reg32 r4349 (rst, clk, in, r4349_out);
	reg32 r4350 (rst, clk, in, r4350_out);
	reg32 r4351 (rst, clk, in, r4351_out);
	reg32 r4352 (rst, clk, in, r4352_out);
	reg32 r4353 (rst, clk, in, r4353_out);
	reg32 r4354 (rst, clk, in, r4354_out);
	reg32 r4355 (rst, clk, in, r4355_out);
	reg32 r4356 (rst, clk, in, r4356_out);
	reg32 r4357 (rst, clk, in, r4357_out);
	reg32 r4358 (rst, clk, in, r4358_out);
	reg32 r4359 (rst, clk, in, r4359_out);
	reg32 r4360 (rst, clk, in, r4360_out);
	reg32 r4361 (rst, clk, in, r4361_out);
	reg32 r4362 (rst, clk, in, r4362_out);
	reg32 r4363 (rst, clk, in, r4363_out);
	reg32 r4364 (rst, clk, in, r4364_out);
	reg32 r4365 (rst, clk, in, r4365_out);
	reg32 r4366 (rst, clk, in, r4366_out);
	reg32 r4367 (rst, clk, in, r4367_out);
	reg32 r4368 (rst, clk, in, r4368_out);
	reg32 r4369 (rst, clk, in, r4369_out);
	reg32 r4370 (rst, clk, in, r4370_out);
	reg32 r4371 (rst, clk, in, r4371_out);
	reg32 r4372 (rst, clk, in, r4372_out);
	reg32 r4373 (rst, clk, in, r4373_out);
	reg32 r4374 (rst, clk, in, r4374_out);
	reg32 r4375 (rst, clk, in, r4375_out);
	reg32 r4376 (rst, clk, in, r4376_out);
	reg32 r4377 (rst, clk, in, r4377_out);
	reg32 r4378 (rst, clk, in, r4378_out);
	reg32 r4379 (rst, clk, in, r4379_out);
	reg32 r4380 (rst, clk, in, r4380_out);
	reg32 r4381 (rst, clk, in, r4381_out);
	reg32 r4382 (rst, clk, in, r4382_out);
	reg32 r4383 (rst, clk, in, r4383_out);
	reg32 r4384 (rst, clk, in, r4384_out);
	reg32 r4385 (rst, clk, in, r4385_out);
	reg32 r4386 (rst, clk, in, r4386_out);
	reg32 r4387 (rst, clk, in, r4387_out);
	reg32 r4388 (rst, clk, in, r4388_out);
	reg32 r4389 (rst, clk, in, r4389_out);
	reg32 r4390 (rst, clk, in, r4390_out);
	reg32 r4391 (rst, clk, in, r4391_out);
	reg32 r4392 (rst, clk, in, r4392_out);
	reg32 r4393 (rst, clk, in, r4393_out);
	reg32 r4394 (rst, clk, in, r4394_out);
	reg32 r4395 (rst, clk, in, r4395_out);
	reg32 r4396 (rst, clk, in, r4396_out);
	reg32 r4397 (rst, clk, in, r4397_out);
	reg32 r4398 (rst, clk, in, r4398_out);
	reg32 r4399 (rst, clk, in, r4399_out);
	reg32 r4400 (rst, clk, in, r4400_out);
	reg32 r4401 (rst, clk, in, r4401_out);
	reg32 r4402 (rst, clk, in, r4402_out);
	reg32 r4403 (rst, clk, in, r4403_out);
	reg32 r4404 (rst, clk, in, r4404_out);
	reg32 r4405 (rst, clk, in, r4405_out);
	reg32 r4406 (rst, clk, in, r4406_out);
	reg32 r4407 (rst, clk, in, r4407_out);
	reg32 r4408 (rst, clk, in, r4408_out);
	reg32 r4409 (rst, clk, in, r4409_out);
	reg32 r4410 (rst, clk, in, r4410_out);
	reg32 r4411 (rst, clk, in, r4411_out);
	reg32 r4412 (rst, clk, in, r4412_out);
	reg32 r4413 (rst, clk, in, r4413_out);
	reg32 r4414 (rst, clk, in, r4414_out);
	reg32 r4415 (rst, clk, in, r4415_out);
	reg32 r4416 (rst, clk, in, r4416_out);
	reg32 r4417 (rst, clk, in, r4417_out);
	reg32 r4418 (rst, clk, in, r4418_out);
	reg32 r4419 (rst, clk, in, r4419_out);
	reg32 r4420 (rst, clk, in, r4420_out);
	reg32 r4421 (rst, clk, in, r4421_out);
	reg32 r4422 (rst, clk, in, r4422_out);
	reg32 r4423 (rst, clk, in, r4423_out);
	reg32 r4424 (rst, clk, in, r4424_out);
	reg32 r4425 (rst, clk, in, r4425_out);
	reg32 r4426 (rst, clk, in, r4426_out);
	reg32 r4427 (rst, clk, in, r4427_out);
	reg32 r4428 (rst, clk, in, r4428_out);
	reg32 r4429 (rst, clk, in, r4429_out);
	reg32 r4430 (rst, clk, in, r4430_out);
	reg32 r4431 (rst, clk, in, r4431_out);
	reg32 r4432 (rst, clk, in, r4432_out);
	reg32 r4433 (rst, clk, in, r4433_out);
	reg32 r4434 (rst, clk, in, r4434_out);
	reg32 r4435 (rst, clk, in, r4435_out);
	reg32 r4436 (rst, clk, in, r4436_out);
	reg32 r4437 (rst, clk, in, r4437_out);
	reg32 r4438 (rst, clk, in, r4438_out);
	reg32 r4439 (rst, clk, in, r4439_out);
	reg32 r4440 (rst, clk, in, r4440_out);
	reg32 r4441 (rst, clk, in, r4441_out);
	reg32 r4442 (rst, clk, in, r4442_out);
	reg32 r4443 (rst, clk, in, r4443_out);
	reg32 r4444 (rst, clk, in, r4444_out);
	reg32 r4445 (rst, clk, in, r4445_out);
	reg32 r4446 (rst, clk, in, r4446_out);
	reg32 r4447 (rst, clk, in, r4447_out);
	reg32 r4448 (rst, clk, in, r4448_out);
	reg32 r4449 (rst, clk, in, r4449_out);
	reg32 r4450 (rst, clk, in, r4450_out);
	reg32 r4451 (rst, clk, in, r4451_out);
	reg32 r4452 (rst, clk, in, r4452_out);
	reg32 r4453 (rst, clk, in, r4453_out);
	reg32 r4454 (rst, clk, in, r4454_out);
	reg32 r4455 (rst, clk, in, r4455_out);
	reg32 r4456 (rst, clk, in, r4456_out);
	reg32 r4457 (rst, clk, in, r4457_out);
	reg32 r4458 (rst, clk, in, r4458_out);
	reg32 r4459 (rst, clk, in, r4459_out);
	reg32 r4460 (rst, clk, in, r4460_out);
	reg32 r4461 (rst, clk, in, r4461_out);
	reg32 r4462 (rst, clk, in, r4462_out);
	reg32 r4463 (rst, clk, in, r4463_out);
	reg32 r4464 (rst, clk, in, r4464_out);
	reg32 r4465 (rst, clk, in, r4465_out);
	reg32 r4466 (rst, clk, in, r4466_out);
	reg32 r4467 (rst, clk, in, r4467_out);
	reg32 r4468 (rst, clk, in, r4468_out);
	reg32 r4469 (rst, clk, in, r4469_out);
	reg32 r4470 (rst, clk, in, r4470_out);
	reg32 r4471 (rst, clk, in, r4471_out);
	reg32 r4472 (rst, clk, in, r4472_out);
	reg32 r4473 (rst, clk, in, r4473_out);
	reg32 r4474 (rst, clk, in, r4474_out);
	reg32 r4475 (rst, clk, in, r4475_out);
	reg32 r4476 (rst, clk, in, r4476_out);
	reg32 r4477 (rst, clk, in, r4477_out);
	reg32 r4478 (rst, clk, in, r4478_out);
	reg32 r4479 (rst, clk, in, r4479_out);
	reg32 r4480 (rst, clk, in, r4480_out);
	reg32 r4481 (rst, clk, in, r4481_out);
	reg32 r4482 (rst, clk, in, r4482_out);
	reg32 r4483 (rst, clk, in, r4483_out);
	reg32 r4484 (rst, clk, in, r4484_out);
	reg32 r4485 (rst, clk, in, r4485_out);
	reg32 r4486 (rst, clk, in, r4486_out);
	reg32 r4487 (rst, clk, in, r4487_out);
	reg32 r4488 (rst, clk, in, r4488_out);
	reg32 r4489 (rst, clk, in, r4489_out);
	reg32 r4490 (rst, clk, in, r4490_out);
	reg32 r4491 (rst, clk, in, r4491_out);
	reg32 r4492 (rst, clk, in, r4492_out);
	reg32 r4493 (rst, clk, in, r4493_out);
	reg32 r4494 (rst, clk, in, r4494_out);
	reg32 r4495 (rst, clk, in, r4495_out);
	reg32 r4496 (rst, clk, in, r4496_out);
	reg32 r4497 (rst, clk, in, r4497_out);
	reg32 r4498 (rst, clk, in, r4498_out);
	reg32 r4499 (rst, clk, in, r4499_out);
	reg32 r4500 (rst, clk, in, r4500_out);
	reg32 r4501 (rst, clk, in, r4501_out);
	reg32 r4502 (rst, clk, in, r4502_out);
	reg32 r4503 (rst, clk, in, r4503_out);
	reg32 r4504 (rst, clk, in, r4504_out);
	reg32 r4505 (rst, clk, in, r4505_out);
	reg32 r4506 (rst, clk, in, r4506_out);
	reg32 r4507 (rst, clk, in, r4507_out);
	reg32 r4508 (rst, clk, in, r4508_out);
	reg32 r4509 (rst, clk, in, r4509_out);
	reg32 r4510 (rst, clk, in, r4510_out);
	reg32 r4511 (rst, clk, in, r4511_out);
	reg32 r4512 (rst, clk, in, r4512_out);
	reg32 r4513 (rst, clk, in, r4513_out);
	reg32 r4514 (rst, clk, in, r4514_out);
	reg32 r4515 (rst, clk, in, r4515_out);
	reg32 r4516 (rst, clk, in, r4516_out);
	reg32 r4517 (rst, clk, in, r4517_out);
	reg32 r4518 (rst, clk, in, r4518_out);
	reg32 r4519 (rst, clk, in, r4519_out);
	reg32 r4520 (rst, clk, in, r4520_out);
	reg32 r4521 (rst, clk, in, r4521_out);
	reg32 r4522 (rst, clk, in, r4522_out);
	reg32 r4523 (rst, clk, in, r4523_out);
	reg32 r4524 (rst, clk, in, r4524_out);
	reg32 r4525 (rst, clk, in, r4525_out);
	reg32 r4526 (rst, clk, in, r4526_out);
	reg32 r4527 (rst, clk, in, r4527_out);
	reg32 r4528 (rst, clk, in, r4528_out);
	reg32 r4529 (rst, clk, in, r4529_out);
	reg32 r4530 (rst, clk, in, r4530_out);
	reg32 r4531 (rst, clk, in, r4531_out);
	reg32 r4532 (rst, clk, in, r4532_out);
	reg32 r4533 (rst, clk, in, r4533_out);
	reg32 r4534 (rst, clk, in, r4534_out);
	reg32 r4535 (rst, clk, in, r4535_out);
	reg32 r4536 (rst, clk, in, r4536_out);
	reg32 r4537 (rst, clk, in, r4537_out);
	reg32 r4538 (rst, clk, in, r4538_out);
	reg32 r4539 (rst, clk, in, r4539_out);
	reg32 r4540 (rst, clk, in, r4540_out);
	reg32 r4541 (rst, clk, in, r4541_out);
	reg32 r4542 (rst, clk, in, r4542_out);
	reg32 r4543 (rst, clk, in, r4543_out);
	reg32 r4544 (rst, clk, in, r4544_out);
	reg32 r4545 (rst, clk, in, r4545_out);
	reg32 r4546 (rst, clk, in, r4546_out);
	reg32 r4547 (rst, clk, in, r4547_out);
	reg32 r4548 (rst, clk, in, r4548_out);
	reg32 r4549 (rst, clk, in, r4549_out);
	reg32 r4550 (rst, clk, in, r4550_out);
	reg32 r4551 (rst, clk, in, r4551_out);
	reg32 r4552 (rst, clk, in, r4552_out);
	reg32 r4553 (rst, clk, in, r4553_out);
	reg32 r4554 (rst, clk, in, r4554_out);
	reg32 r4555 (rst, clk, in, r4555_out);
	reg32 r4556 (rst, clk, in, r4556_out);
	reg32 r4557 (rst, clk, in, r4557_out);
	reg32 r4558 (rst, clk, in, r4558_out);
	reg32 r4559 (rst, clk, in, r4559_out);
	reg32 r4560 (rst, clk, in, r4560_out);
	reg32 r4561 (rst, clk, in, r4561_out);
	reg32 r4562 (rst, clk, in, r4562_out);
	reg32 r4563 (rst, clk, in, r4563_out);
	reg32 r4564 (rst, clk, in, r4564_out);
	reg32 r4565 (rst, clk, in, r4565_out);
	reg32 r4566 (rst, clk, in, r4566_out);
	reg32 r4567 (rst, clk, in, r4567_out);
	reg32 r4568 (rst, clk, in, r4568_out);
	reg32 r4569 (rst, clk, in, r4569_out);
	reg32 r4570 (rst, clk, in, r4570_out);
	reg32 r4571 (rst, clk, in, r4571_out);
	reg32 r4572 (rst, clk, in, r4572_out);
	reg32 r4573 (rst, clk, in, r4573_out);
	reg32 r4574 (rst, clk, in, r4574_out);
	reg32 r4575 (rst, clk, in, r4575_out);
	reg32 r4576 (rst, clk, in, r4576_out);
	reg32 r4577 (rst, clk, in, r4577_out);
	reg32 r4578 (rst, clk, in, r4578_out);
	reg32 r4579 (rst, clk, in, r4579_out);
	reg32 r4580 (rst, clk, in, r4580_out);
	reg32 r4581 (rst, clk, in, r4581_out);
	reg32 r4582 (rst, clk, in, r4582_out);
	reg32 r4583 (rst, clk, in, r4583_out);
	reg32 r4584 (rst, clk, in, r4584_out);
	reg32 r4585 (rst, clk, in, r4585_out);
	reg32 r4586 (rst, clk, in, r4586_out);
	reg32 r4587 (rst, clk, in, r4587_out);
	reg32 r4588 (rst, clk, in, r4588_out);
	reg32 r4589 (rst, clk, in, r4589_out);
	reg32 r4590 (rst, clk, in, r4590_out);
	reg32 r4591 (rst, clk, in, r4591_out);
	reg32 r4592 (rst, clk, in, r4592_out);
	reg32 r4593 (rst, clk, in, r4593_out);
	reg32 r4594 (rst, clk, in, r4594_out);
	reg32 r4595 (rst, clk, in, r4595_out);
	reg32 r4596 (rst, clk, in, r4596_out);
	reg32 r4597 (rst, clk, in, r4597_out);
	reg32 r4598 (rst, clk, in, r4598_out);
	reg32 r4599 (rst, clk, in, r4599_out);
	reg32 r4600 (rst, clk, in, r4600_out);
	reg32 r4601 (rst, clk, in, r4601_out);
	reg32 r4602 (rst, clk, in, r4602_out);
	reg32 r4603 (rst, clk, in, r4603_out);
	reg32 r4604 (rst, clk, in, r4604_out);
	reg32 r4605 (rst, clk, in, r4605_out);
	reg32 r4606 (rst, clk, in, r4606_out);
	reg32 r4607 (rst, clk, in, r4607_out);
	reg32 r4608 (rst, clk, in, r4608_out);
	reg32 r4609 (rst, clk, in, r4609_out);
	reg32 r4610 (rst, clk, in, r4610_out);
	reg32 r4611 (rst, clk, in, r4611_out);
	reg32 r4612 (rst, clk, in, r4612_out);
	reg32 r4613 (rst, clk, in, r4613_out);
	reg32 r4614 (rst, clk, in, r4614_out);
	reg32 r4615 (rst, clk, in, r4615_out);
	reg32 r4616 (rst, clk, in, r4616_out);
	reg32 r4617 (rst, clk, in, r4617_out);
	reg32 r4618 (rst, clk, in, r4618_out);
	reg32 r4619 (rst, clk, in, r4619_out);
	reg32 r4620 (rst, clk, in, r4620_out);
	reg32 r4621 (rst, clk, in, r4621_out);
	reg32 r4622 (rst, clk, in, r4622_out);
	reg32 r4623 (rst, clk, in, r4623_out);
	reg32 r4624 (rst, clk, in, r4624_out);
	reg32 r4625 (rst, clk, in, r4625_out);
	reg32 r4626 (rst, clk, in, r4626_out);
	reg32 r4627 (rst, clk, in, r4627_out);
	reg32 r4628 (rst, clk, in, r4628_out);
	reg32 r4629 (rst, clk, in, r4629_out);
	reg32 r4630 (rst, clk, in, r4630_out);
	reg32 r4631 (rst, clk, in, r4631_out);
	reg32 r4632 (rst, clk, in, r4632_out);
	reg32 r4633 (rst, clk, in, r4633_out);
	reg32 r4634 (rst, clk, in, r4634_out);
	reg32 r4635 (rst, clk, in, r4635_out);
	reg32 r4636 (rst, clk, in, r4636_out);
	reg32 r4637 (rst, clk, in, r4637_out);
	reg32 r4638 (rst, clk, in, r4638_out);
	reg32 r4639 (rst, clk, in, r4639_out);
	reg32 r4640 (rst, clk, in, r4640_out);
	reg32 r4641 (rst, clk, in, r4641_out);
	reg32 r4642 (rst, clk, in, r4642_out);
	reg32 r4643 (rst, clk, in, r4643_out);
	reg32 r4644 (rst, clk, in, r4644_out);
	reg32 r4645 (rst, clk, in, r4645_out);
	reg32 r4646 (rst, clk, in, r4646_out);
	reg32 r4647 (rst, clk, in, r4647_out);
	reg32 r4648 (rst, clk, in, r4648_out);
	reg32 r4649 (rst, clk, in, r4649_out);
	reg32 r4650 (rst, clk, in, r4650_out);
	reg32 r4651 (rst, clk, in, r4651_out);
	reg32 r4652 (rst, clk, in, r4652_out);
	reg32 r4653 (rst, clk, in, r4653_out);
	reg32 r4654 (rst, clk, in, r4654_out);
	reg32 r4655 (rst, clk, in, r4655_out);
	reg32 r4656 (rst, clk, in, r4656_out);
	reg32 r4657 (rst, clk, in, r4657_out);
	reg32 r4658 (rst, clk, in, r4658_out);
	reg32 r4659 (rst, clk, in, r4659_out);
	reg32 r4660 (rst, clk, in, r4660_out);
	reg32 r4661 (rst, clk, in, r4661_out);
	reg32 r4662 (rst, clk, in, r4662_out);
	reg32 r4663 (rst, clk, in, r4663_out);
	reg32 r4664 (rst, clk, in, r4664_out);
	reg32 r4665 (rst, clk, in, r4665_out);
	reg32 r4666 (rst, clk, in, r4666_out);
	reg32 r4667 (rst, clk, in, r4667_out);
	reg32 r4668 (rst, clk, in, r4668_out);
	reg32 r4669 (rst, clk, in, r4669_out);
	reg32 r4670 (rst, clk, in, r4670_out);
	reg32 r4671 (rst, clk, in, r4671_out);
	reg32 r4672 (rst, clk, in, r4672_out);
	reg32 r4673 (rst, clk, in, r4673_out);
	reg32 r4674 (rst, clk, in, r4674_out);
	reg32 r4675 (rst, clk, in, r4675_out);
	reg32 r4676 (rst, clk, in, r4676_out);
	reg32 r4677 (rst, clk, in, r4677_out);
	reg32 r4678 (rst, clk, in, r4678_out);
	reg32 r4679 (rst, clk, in, r4679_out);
	reg32 r4680 (rst, clk, in, r4680_out);
	reg32 r4681 (rst, clk, in, r4681_out);
	reg32 r4682 (rst, clk, in, r4682_out);
	reg32 r4683 (rst, clk, in, r4683_out);
	reg32 r4684 (rst, clk, in, r4684_out);
	reg32 r4685 (rst, clk, in, r4685_out);
	reg32 r4686 (rst, clk, in, r4686_out);
	reg32 r4687 (rst, clk, in, r4687_out);
	reg32 r4688 (rst, clk, in, r4688_out);
	reg32 r4689 (rst, clk, in, r4689_out);
	reg32 r4690 (rst, clk, in, r4690_out);
	reg32 r4691 (rst, clk, in, r4691_out);
	reg32 r4692 (rst, clk, in, r4692_out);
	reg32 r4693 (rst, clk, in, r4693_out);
	reg32 r4694 (rst, clk, in, r4694_out);
	reg32 r4695 (rst, clk, in, r4695_out);
	reg32 r4696 (rst, clk, in, r4696_out);
	reg32 r4697 (rst, clk, in, r4697_out);
	reg32 r4698 (rst, clk, in, r4698_out);
	reg32 r4699 (rst, clk, in, r4699_out);
	reg32 r4700 (rst, clk, in, r4700_out);
	reg32 r4701 (rst, clk, in, r4701_out);
	reg32 r4702 (rst, clk, in, r4702_out);
	reg32 r4703 (rst, clk, in, r4703_out);
	reg32 r4704 (rst, clk, in, r4704_out);
	reg32 r4705 (rst, clk, in, r4705_out);
	reg32 r4706 (rst, clk, in, r4706_out);
	reg32 r4707 (rst, clk, in, r4707_out);
	reg32 r4708 (rst, clk, in, r4708_out);
	reg32 r4709 (rst, clk, in, r4709_out);
	reg32 r4710 (rst, clk, in, r4710_out);
	reg32 r4711 (rst, clk, in, r4711_out);
	reg32 r4712 (rst, clk, in, r4712_out);
	reg32 r4713 (rst, clk, in, r4713_out);
	reg32 r4714 (rst, clk, in, r4714_out);
	reg32 r4715 (rst, clk, in, r4715_out);
	reg32 r4716 (rst, clk, in, r4716_out);
	reg32 r4717 (rst, clk, in, r4717_out);
	reg32 r4718 (rst, clk, in, r4718_out);
	reg32 r4719 (rst, clk, in, r4719_out);
	reg32 r4720 (rst, clk, in, r4720_out);
	reg32 r4721 (rst, clk, in, r4721_out);
	reg32 r4722 (rst, clk, in, r4722_out);
	reg32 r4723 (rst, clk, in, r4723_out);
	reg32 r4724 (rst, clk, in, r4724_out);
	reg32 r4725 (rst, clk, in, r4725_out);
	reg32 r4726 (rst, clk, in, r4726_out);
	reg32 r4727 (rst, clk, in, r4727_out);
	reg32 r4728 (rst, clk, in, r4728_out);
	reg32 r4729 (rst, clk, in, r4729_out);
	reg32 r4730 (rst, clk, in, r4730_out);
	reg32 r4731 (rst, clk, in, r4731_out);
	reg32 r4732 (rst, clk, in, r4732_out);
	reg32 r4733 (rst, clk, in, r4733_out);
	reg32 r4734 (rst, clk, in, r4734_out);
	reg32 r4735 (rst, clk, in, r4735_out);
	reg32 r4736 (rst, clk, in, r4736_out);
	reg32 r4737 (rst, clk, in, r4737_out);
	reg32 r4738 (rst, clk, in, r4738_out);
	reg32 r4739 (rst, clk, in, r4739_out);
	reg32 r4740 (rst, clk, in, r4740_out);
	reg32 r4741 (rst, clk, in, r4741_out);
	reg32 r4742 (rst, clk, in, r4742_out);
	reg32 r4743 (rst, clk, in, r4743_out);
	reg32 r4744 (rst, clk, in, r4744_out);
	reg32 r4745 (rst, clk, in, r4745_out);
	reg32 r4746 (rst, clk, in, r4746_out);
	reg32 r4747 (rst, clk, in, r4747_out);
	reg32 r4748 (rst, clk, in, r4748_out);
	reg32 r4749 (rst, clk, in, r4749_out);
	reg32 r4750 (rst, clk, in, r4750_out);
	reg32 r4751 (rst, clk, in, r4751_out);
	reg32 r4752 (rst, clk, in, r4752_out);
	reg32 r4753 (rst, clk, in, r4753_out);
	reg32 r4754 (rst, clk, in, r4754_out);
	reg32 r4755 (rst, clk, in, r4755_out);
	reg32 r4756 (rst, clk, in, r4756_out);
	reg32 r4757 (rst, clk, in, r4757_out);
	reg32 r4758 (rst, clk, in, r4758_out);
	reg32 r4759 (rst, clk, in, r4759_out);
	reg32 r4760 (rst, clk, in, r4760_out);
	reg32 r4761 (rst, clk, in, r4761_out);
	reg32 r4762 (rst, clk, in, r4762_out);
	reg32 r4763 (rst, clk, in, r4763_out);
	reg32 r4764 (rst, clk, in, r4764_out);
	reg32 r4765 (rst, clk, in, r4765_out);
	reg32 r4766 (rst, clk, in, r4766_out);
	reg32 r4767 (rst, clk, in, r4767_out);
	reg32 r4768 (rst, clk, in, r4768_out);
	reg32 r4769 (rst, clk, in, r4769_out);
	reg32 r4770 (rst, clk, in, r4770_out);
	reg32 r4771 (rst, clk, in, r4771_out);
	reg32 r4772 (rst, clk, in, r4772_out);
	reg32 r4773 (rst, clk, in, r4773_out);
	reg32 r4774 (rst, clk, in, r4774_out);
	reg32 r4775 (rst, clk, in, r4775_out);
	reg32 r4776 (rst, clk, in, r4776_out);
	reg32 r4777 (rst, clk, in, r4777_out);
	reg32 r4778 (rst, clk, in, r4778_out);
	reg32 r4779 (rst, clk, in, r4779_out);
	reg32 r4780 (rst, clk, in, r4780_out);
	reg32 r4781 (rst, clk, in, r4781_out);
	reg32 r4782 (rst, clk, in, r4782_out);
	reg32 r4783 (rst, clk, in, r4783_out);
	reg32 r4784 (rst, clk, in, r4784_out);
	reg32 r4785 (rst, clk, in, r4785_out);
	reg32 r4786 (rst, clk, in, r4786_out);
	reg32 r4787 (rst, clk, in, r4787_out);
	reg32 r4788 (rst, clk, in, r4788_out);
	reg32 r4789 (rst, clk, in, r4789_out);
	reg32 r4790 (rst, clk, in, r4790_out);
	reg32 r4791 (rst, clk, in, r4791_out);
	reg32 r4792 (rst, clk, in, r4792_out);
	reg32 r4793 (rst, clk, in, r4793_out);
	reg32 r4794 (rst, clk, in, r4794_out);
	reg32 r4795 (rst, clk, in, r4795_out);
	reg32 r4796 (rst, clk, in, r4796_out);
	reg32 r4797 (rst, clk, in, r4797_out);
	reg32 r4798 (rst, clk, in, r4798_out);
	reg32 r4799 (rst, clk, in, r4799_out);
	reg32 r4800 (rst, clk, in, r4800_out);
	reg32 r4801 (rst, clk, in, r4801_out);
	reg32 r4802 (rst, clk, in, r4802_out);
	reg32 r4803 (rst, clk, in, r4803_out);
	reg32 r4804 (rst, clk, in, r4804_out);
	reg32 r4805 (rst, clk, in, r4805_out);
	reg32 r4806 (rst, clk, in, r4806_out);
	reg32 r4807 (rst, clk, in, r4807_out);
	reg32 r4808 (rst, clk, in, r4808_out);
	reg32 r4809 (rst, clk, in, r4809_out);
	reg32 r4810 (rst, clk, in, r4810_out);
	reg32 r4811 (rst, clk, in, r4811_out);
	reg32 r4812 (rst, clk, in, r4812_out);
	reg32 r4813 (rst, clk, in, r4813_out);
	reg32 r4814 (rst, clk, in, r4814_out);
	reg32 r4815 (rst, clk, in, r4815_out);
	reg32 r4816 (rst, clk, in, r4816_out);
	reg32 r4817 (rst, clk, in, r4817_out);
	reg32 r4818 (rst, clk, in, r4818_out);
	reg32 r4819 (rst, clk, in, r4819_out);
	reg32 r4820 (rst, clk, in, r4820_out);
	reg32 r4821 (rst, clk, in, r4821_out);
	reg32 r4822 (rst, clk, in, r4822_out);
	reg32 r4823 (rst, clk, in, r4823_out);
	reg32 r4824 (rst, clk, in, r4824_out);
	reg32 r4825 (rst, clk, in, r4825_out);
	reg32 r4826 (rst, clk, in, r4826_out);
	reg32 r4827 (rst, clk, in, r4827_out);
	reg32 r4828 (rst, clk, in, r4828_out);
	reg32 r4829 (rst, clk, in, r4829_out);
	reg32 r4830 (rst, clk, in, r4830_out);
	reg32 r4831 (rst, clk, in, r4831_out);
	reg32 r4832 (rst, clk, in, r4832_out);
	reg32 r4833 (rst, clk, in, r4833_out);
	reg32 r4834 (rst, clk, in, r4834_out);
	reg32 r4835 (rst, clk, in, r4835_out);
	reg32 r4836 (rst, clk, in, r4836_out);
	reg32 r4837 (rst, clk, in, r4837_out);
	reg32 r4838 (rst, clk, in, r4838_out);
	reg32 r4839 (rst, clk, in, r4839_out);
	reg32 r4840 (rst, clk, in, r4840_out);
	reg32 r4841 (rst, clk, in, r4841_out);
	reg32 r4842 (rst, clk, in, r4842_out);
	reg32 r4843 (rst, clk, in, r4843_out);
	reg32 r4844 (rst, clk, in, r4844_out);
	reg32 r4845 (rst, clk, in, r4845_out);
	reg32 r4846 (rst, clk, in, r4846_out);
	reg32 r4847 (rst, clk, in, r4847_out);
	reg32 r4848 (rst, clk, in, r4848_out);
	reg32 r4849 (rst, clk, in, r4849_out);
	reg32 r4850 (rst, clk, in, r4850_out);
	reg32 r4851 (rst, clk, in, r4851_out);
	reg32 r4852 (rst, clk, in, r4852_out);
	reg32 r4853 (rst, clk, in, r4853_out);
	reg32 r4854 (rst, clk, in, r4854_out);
	reg32 r4855 (rst, clk, in, r4855_out);
	reg32 r4856 (rst, clk, in, r4856_out);
	reg32 r4857 (rst, clk, in, r4857_out);
	reg32 r4858 (rst, clk, in, r4858_out);
	reg32 r4859 (rst, clk, in, r4859_out);
	reg32 r4860 (rst, clk, in, r4860_out);
	reg32 r4861 (rst, clk, in, r4861_out);
	reg32 r4862 (rst, clk, in, r4862_out);
	reg32 r4863 (rst, clk, in, r4863_out);
	reg32 r4864 (rst, clk, in, r4864_out);
	reg32 r4865 (rst, clk, in, r4865_out);
	reg32 r4866 (rst, clk, in, r4866_out);
	reg32 r4867 (rst, clk, in, r4867_out);
	reg32 r4868 (rst, clk, in, r4868_out);
	reg32 r4869 (rst, clk, in, r4869_out);
	reg32 r4870 (rst, clk, in, r4870_out);
	reg32 r4871 (rst, clk, in, r4871_out);
	reg32 r4872 (rst, clk, in, r4872_out);
	reg32 r4873 (rst, clk, in, r4873_out);
	reg32 r4874 (rst, clk, in, r4874_out);
	reg32 r4875 (rst, clk, in, r4875_out);
	reg32 r4876 (rst, clk, in, r4876_out);
	reg32 r4877 (rst, clk, in, r4877_out);
	reg32 r4878 (rst, clk, in, r4878_out);
	reg32 r4879 (rst, clk, in, r4879_out);
	reg32 r4880 (rst, clk, in, r4880_out);
	reg32 r4881 (rst, clk, in, r4881_out);
	reg32 r4882 (rst, clk, in, r4882_out);
	reg32 r4883 (rst, clk, in, r4883_out);
	reg32 r4884 (rst, clk, in, r4884_out);
	reg32 r4885 (rst, clk, in, r4885_out);
	reg32 r4886 (rst, clk, in, r4886_out);
	reg32 r4887 (rst, clk, in, r4887_out);
	reg32 r4888 (rst, clk, in, r4888_out);
	reg32 r4889 (rst, clk, in, r4889_out);
	reg32 r4890 (rst, clk, in, r4890_out);
	reg32 r4891 (rst, clk, in, r4891_out);
	reg32 r4892 (rst, clk, in, r4892_out);
	reg32 r4893 (rst, clk, in, r4893_out);
	reg32 r4894 (rst, clk, in, r4894_out);
	reg32 r4895 (rst, clk, in, r4895_out);
	reg32 r4896 (rst, clk, in, r4896_out);
	reg32 r4897 (rst, clk, in, r4897_out);
	reg32 r4898 (rst, clk, in, r4898_out);
	reg32 r4899 (rst, clk, in, r4899_out);
	reg32 r4900 (rst, clk, in, r4900_out);
	reg32 r4901 (rst, clk, in, r4901_out);
	reg32 r4902 (rst, clk, in, r4902_out);
	reg32 r4903 (rst, clk, in, r4903_out);
	reg32 r4904 (rst, clk, in, r4904_out);
	reg32 r4905 (rst, clk, in, r4905_out);
	reg32 r4906 (rst, clk, in, r4906_out);
	reg32 r4907 (rst, clk, in, r4907_out);
	reg32 r4908 (rst, clk, in, r4908_out);
	reg32 r4909 (rst, clk, in, r4909_out);
	reg32 r4910 (rst, clk, in, r4910_out);
	reg32 r4911 (rst, clk, in, r4911_out);
	reg32 r4912 (rst, clk, in, r4912_out);
	reg32 r4913 (rst, clk, in, r4913_out);
	reg32 r4914 (rst, clk, in, r4914_out);
	reg32 r4915 (rst, clk, in, r4915_out);
	reg32 r4916 (rst, clk, in, r4916_out);
	reg32 r4917 (rst, clk, in, r4917_out);
	reg32 r4918 (rst, clk, in, r4918_out);
	reg32 r4919 (rst, clk, in, r4919_out);
	reg32 r4920 (rst, clk, in, r4920_out);
	reg32 r4921 (rst, clk, in, r4921_out);
	reg32 r4922 (rst, clk, in, r4922_out);
	reg32 r4923 (rst, clk, in, r4923_out);
	reg32 r4924 (rst, clk, in, r4924_out);
	reg32 r4925 (rst, clk, in, r4925_out);
	reg32 r4926 (rst, clk, in, r4926_out);
	reg32 r4927 (rst, clk, in, r4927_out);
	reg32 r4928 (rst, clk, in, r4928_out);
	reg32 r4929 (rst, clk, in, r4929_out);
	reg32 r4930 (rst, clk, in, r4930_out);
	reg32 r4931 (rst, clk, in, r4931_out);
	reg32 r4932 (rst, clk, in, r4932_out);
	reg32 r4933 (rst, clk, in, r4933_out);
	reg32 r4934 (rst, clk, in, r4934_out);
	reg32 r4935 (rst, clk, in, r4935_out);
	reg32 r4936 (rst, clk, in, r4936_out);
	reg32 r4937 (rst, clk, in, r4937_out);
	reg32 r4938 (rst, clk, in, r4938_out);
	reg32 r4939 (rst, clk, in, r4939_out);
	reg32 r4940 (rst, clk, in, r4940_out);
	reg32 r4941 (rst, clk, in, r4941_out);
	reg32 r4942 (rst, clk, in, r4942_out);
	reg32 r4943 (rst, clk, in, r4943_out);
	reg32 r4944 (rst, clk, in, r4944_out);
	reg32 r4945 (rst, clk, in, r4945_out);
	reg32 r4946 (rst, clk, in, r4946_out);
	reg32 r4947 (rst, clk, in, r4947_out);
	reg32 r4948 (rst, clk, in, r4948_out);
	reg32 r4949 (rst, clk, in, r4949_out);
	reg32 r4950 (rst, clk, in, r4950_out);
	reg32 r4951 (rst, clk, in, r4951_out);
	reg32 r4952 (rst, clk, in, r4952_out);
	reg32 r4953 (rst, clk, in, r4953_out);
	reg32 r4954 (rst, clk, in, r4954_out);
	reg32 r4955 (rst, clk, in, r4955_out);
	reg32 r4956 (rst, clk, in, r4956_out);
	reg32 r4957 (rst, clk, in, r4957_out);
	reg32 r4958 (rst, clk, in, r4958_out);
	reg32 r4959 (rst, clk, in, r4959_out);
	reg32 r4960 (rst, clk, in, r4960_out);
	reg32 r4961 (rst, clk, in, r4961_out);
	reg32 r4962 (rst, clk, in, r4962_out);
	reg32 r4963 (rst, clk, in, r4963_out);
	reg32 r4964 (rst, clk, in, r4964_out);
	reg32 r4965 (rst, clk, in, r4965_out);
	reg32 r4966 (rst, clk, in, r4966_out);
	reg32 r4967 (rst, clk, in, r4967_out);
	reg32 r4968 (rst, clk, in, r4968_out);
	reg32 r4969 (rst, clk, in, r4969_out);
	reg32 r4970 (rst, clk, in, r4970_out);
	reg32 r4971 (rst, clk, in, r4971_out);
	reg32 r4972 (rst, clk, in, r4972_out);
	reg32 r4973 (rst, clk, in, r4973_out);
	reg32 r4974 (rst, clk, in, r4974_out);
	reg32 r4975 (rst, clk, in, r4975_out);
	reg32 r4976 (rst, clk, in, r4976_out);
	reg32 r4977 (rst, clk, in, r4977_out);
	reg32 r4978 (rst, clk, in, r4978_out);
	reg32 r4979 (rst, clk, in, r4979_out);
	reg32 r4980 (rst, clk, in, r4980_out);
	reg32 r4981 (rst, clk, in, r4981_out);
	reg32 r4982 (rst, clk, in, r4982_out);
	reg32 r4983 (rst, clk, in, r4983_out);
	reg32 r4984 (rst, clk, in, r4984_out);
	reg32 r4985 (rst, clk, in, r4985_out);
	reg32 r4986 (rst, clk, in, r4986_out);
	reg32 r4987 (rst, clk, in, r4987_out);
	reg32 r4988 (rst, clk, in, r4988_out);
	reg32 r4989 (rst, clk, in, r4989_out);
	reg32 r4990 (rst, clk, in, r4990_out);
	reg32 r4991 (rst, clk, in, r4991_out);
	reg32 r4992 (rst, clk, in, r4992_out);
	reg32 r4993 (rst, clk, in, r4993_out);
	reg32 r4994 (rst, clk, in, r4994_out);
	reg32 r4995 (rst, clk, in, r4995_out);
	reg32 r4996 (rst, clk, in, r4996_out);
	reg32 r4997 (rst, clk, in, r4997_out);
	reg32 r4998 (rst, clk, in, r4998_out);
	reg32 r4999 (rst, clk, in, r4999_out);
	reg32 r5000 (rst, clk, in, r5000_out);
	reg32 r5001 (rst, clk, in, r5001_out);
	reg32 r5002 (rst, clk, in, r5002_out);
	reg32 r5003 (rst, clk, in, r5003_out);
	reg32 r5004 (rst, clk, in, r5004_out);
	reg32 r5005 (rst, clk, in, r5005_out);
	reg32 r5006 (rst, clk, in, r5006_out);
	reg32 r5007 (rst, clk, in, r5007_out);
	reg32 r5008 (rst, clk, in, r5008_out);
	reg32 r5009 (rst, clk, in, r5009_out);
	reg32 r5010 (rst, clk, in, r5010_out);
	reg32 r5011 (rst, clk, in, r5011_out);
	reg32 r5012 (rst, clk, in, r5012_out);
	reg32 r5013 (rst, clk, in, r5013_out);
	reg32 r5014 (rst, clk, in, r5014_out);
	reg32 r5015 (rst, clk, in, r5015_out);
	reg32 r5016 (rst, clk, in, r5016_out);
	reg32 r5017 (rst, clk, in, r5017_out);
	reg32 r5018 (rst, clk, in, r5018_out);
	reg32 r5019 (rst, clk, in, r5019_out);
	reg32 r5020 (rst, clk, in, r5020_out);
	reg32 r5021 (rst, clk, in, r5021_out);
	reg32 r5022 (rst, clk, in, r5022_out);
	reg32 r5023 (rst, clk, in, r5023_out);
	reg32 r5024 (rst, clk, in, r5024_out);
	reg32 r5025 (rst, clk, in, r5025_out);
	reg32 r5026 (rst, clk, in, r5026_out);
	reg32 r5027 (rst, clk, in, r5027_out);
	reg32 r5028 (rst, clk, in, r5028_out);
	reg32 r5029 (rst, clk, in, r5029_out);
	reg32 r5030 (rst, clk, in, r5030_out);
	reg32 r5031 (rst, clk, in, r5031_out);
	reg32 r5032 (rst, clk, in, r5032_out);
	reg32 r5033 (rst, clk, in, r5033_out);
	reg32 r5034 (rst, clk, in, r5034_out);
	reg32 r5035 (rst, clk, in, r5035_out);
	reg32 r5036 (rst, clk, in, r5036_out);
	reg32 r5037 (rst, clk, in, r5037_out);
	reg32 r5038 (rst, clk, in, r5038_out);
	reg32 r5039 (rst, clk, in, r5039_out);
	reg32 r5040 (rst, clk, in, r5040_out);
	reg32 r5041 (rst, clk, in, r5041_out);
	reg32 r5042 (rst, clk, in, r5042_out);
	reg32 r5043 (rst, clk, in, r5043_out);
	reg32 r5044 (rst, clk, in, r5044_out);
	reg32 r5045 (rst, clk, in, r5045_out);
	reg32 r5046 (rst, clk, in, r5046_out);
	reg32 r5047 (rst, clk, in, r5047_out);
	reg32 r5048 (rst, clk, in, r5048_out);
	reg32 r5049 (rst, clk, in, r5049_out);
	reg32 r5050 (rst, clk, in, r5050_out);
	reg32 r5051 (rst, clk, in, r5051_out);
	reg32 r5052 (rst, clk, in, r5052_out);
	reg32 r5053 (rst, clk, in, r5053_out);
	reg32 r5054 (rst, clk, in, r5054_out);
	reg32 r5055 (rst, clk, in, r5055_out);
	reg32 r5056 (rst, clk, in, r5056_out);
	reg32 r5057 (rst, clk, in, r5057_out);
	reg32 r5058 (rst, clk, in, r5058_out);
	reg32 r5059 (rst, clk, in, r5059_out);
	reg32 r5060 (rst, clk, in, r5060_out);
	reg32 r5061 (rst, clk, in, r5061_out);
	reg32 r5062 (rst, clk, in, r5062_out);
	reg32 r5063 (rst, clk, in, r5063_out);
	reg32 r5064 (rst, clk, in, r5064_out);
	reg32 r5065 (rst, clk, in, r5065_out);
	reg32 r5066 (rst, clk, in, r5066_out);
	reg32 r5067 (rst, clk, in, r5067_out);
	reg32 r5068 (rst, clk, in, r5068_out);
	reg32 r5069 (rst, clk, in, r5069_out);
	reg32 r5070 (rst, clk, in, r5070_out);
	reg32 r5071 (rst, clk, in, r5071_out);
	reg32 r5072 (rst, clk, in, r5072_out);
	reg32 r5073 (rst, clk, in, r5073_out);
	reg32 r5074 (rst, clk, in, r5074_out);
	reg32 r5075 (rst, clk, in, r5075_out);
	reg32 r5076 (rst, clk, in, r5076_out);
	reg32 r5077 (rst, clk, in, r5077_out);
	reg32 r5078 (rst, clk, in, r5078_out);
	reg32 r5079 (rst, clk, in, r5079_out);
	reg32 r5080 (rst, clk, in, r5080_out);
	reg32 r5081 (rst, clk, in, r5081_out);
	reg32 r5082 (rst, clk, in, r5082_out);
	reg32 r5083 (rst, clk, in, r5083_out);
	reg32 r5084 (rst, clk, in, r5084_out);
	reg32 r5085 (rst, clk, in, r5085_out);
	reg32 r5086 (rst, clk, in, r5086_out);
	reg32 r5087 (rst, clk, in, r5087_out);
	reg32 r5088 (rst, clk, in, r5088_out);
	reg32 r5089 (rst, clk, in, r5089_out);
	reg32 r5090 (rst, clk, in, r5090_out);
	reg32 r5091 (rst, clk, in, r5091_out);
	reg32 r5092 (rst, clk, in, r5092_out);
	reg32 r5093 (rst, clk, in, r5093_out);
	reg32 r5094 (rst, clk, in, r5094_out);
	reg32 r5095 (rst, clk, in, r5095_out);
	reg32 r5096 (rst, clk, in, r5096_out);
	reg32 r5097 (rst, clk, in, r5097_out);
	reg32 r5098 (rst, clk, in, r5098_out);
	reg32 r5099 (rst, clk, in, r5099_out);
	reg32 r5100 (rst, clk, in, r5100_out);
	reg32 r5101 (rst, clk, in, r5101_out);
	reg32 r5102 (rst, clk, in, r5102_out);
	reg32 r5103 (rst, clk, in, r5103_out);
	reg32 r5104 (rst, clk, in, r5104_out);
	reg32 r5105 (rst, clk, in, r5105_out);
	reg32 r5106 (rst, clk, in, r5106_out);
	reg32 r5107 (rst, clk, in, r5107_out);
	reg32 r5108 (rst, clk, in, r5108_out);
	reg32 r5109 (rst, clk, in, r5109_out);
	reg32 r5110 (rst, clk, in, r5110_out);
	reg32 r5111 (rst, clk, in, r5111_out);
	reg32 r5112 (rst, clk, in, r5112_out);
	reg32 r5113 (rst, clk, in, r5113_out);
	reg32 r5114 (rst, clk, in, r5114_out);
	reg32 r5115 (rst, clk, in, r5115_out);
	reg32 r5116 (rst, clk, in, r5116_out);
	reg32 r5117 (rst, clk, in, r5117_out);
	reg32 r5118 (rst, clk, in, r5118_out);
	reg32 r5119 (rst, clk, in, r5119_out);
	reg32 r5120 (rst, clk, in, r5120_out);
	reg32 r5121 (rst, clk, in, r5121_out);
	reg32 r5122 (rst, clk, in, r5122_out);
	reg32 r5123 (rst, clk, in, r5123_out);
	reg32 r5124 (rst, clk, in, r5124_out);
	reg32 r5125 (rst, clk, in, r5125_out);
	reg32 r5126 (rst, clk, in, r5126_out);
	reg32 r5127 (rst, clk, in, r5127_out);
	reg32 r5128 (rst, clk, in, r5128_out);
	reg32 r5129 (rst, clk, in, r5129_out);
	reg32 r5130 (rst, clk, in, r5130_out);
	reg32 r5131 (rst, clk, in, r5131_out);
	reg32 r5132 (rst, clk, in, r5132_out);
	reg32 r5133 (rst, clk, in, r5133_out);
	reg32 r5134 (rst, clk, in, r5134_out);
	reg32 r5135 (rst, clk, in, r5135_out);
	reg32 r5136 (rst, clk, in, r5136_out);
	reg32 r5137 (rst, clk, in, r5137_out);
	reg32 r5138 (rst, clk, in, r5138_out);
	reg32 r5139 (rst, clk, in, r5139_out);
	reg32 r5140 (rst, clk, in, r5140_out);
	reg32 r5141 (rst, clk, in, r5141_out);
	reg32 r5142 (rst, clk, in, r5142_out);
	reg32 r5143 (rst, clk, in, r5143_out);
	reg32 r5144 (rst, clk, in, r5144_out);
	reg32 r5145 (rst, clk, in, r5145_out);
	reg32 r5146 (rst, clk, in, r5146_out);
	reg32 r5147 (rst, clk, in, r5147_out);
	reg32 r5148 (rst, clk, in, r5148_out);
	reg32 r5149 (rst, clk, in, r5149_out);
	reg32 r5150 (rst, clk, in, r5150_out);
	reg32 r5151 (rst, clk, in, r5151_out);
	reg32 r5152 (rst, clk, in, r5152_out);
	reg32 r5153 (rst, clk, in, r5153_out);
	reg32 r5154 (rst, clk, in, r5154_out);
	reg32 r5155 (rst, clk, in, r5155_out);
	reg32 r5156 (rst, clk, in, r5156_out);
	reg32 r5157 (rst, clk, in, r5157_out);
	reg32 r5158 (rst, clk, in, r5158_out);
	reg32 r5159 (rst, clk, in, r5159_out);
	reg32 r5160 (rst, clk, in, r5160_out);
	reg32 r5161 (rst, clk, in, r5161_out);
	reg32 r5162 (rst, clk, in, r5162_out);
	reg32 r5163 (rst, clk, in, r5163_out);
	reg32 r5164 (rst, clk, in, r5164_out);
	reg32 r5165 (rst, clk, in, r5165_out);
	reg32 r5166 (rst, clk, in, r5166_out);
	reg32 r5167 (rst, clk, in, r5167_out);
	reg32 r5168 (rst, clk, in, r5168_out);
	reg32 r5169 (rst, clk, in, r5169_out);
	reg32 r5170 (rst, clk, in, r5170_out);
	reg32 r5171 (rst, clk, in, r5171_out);
	reg32 r5172 (rst, clk, in, r5172_out);
	reg32 r5173 (rst, clk, in, r5173_out);
	reg32 r5174 (rst, clk, in, r5174_out);
	reg32 r5175 (rst, clk, in, r5175_out);
	reg32 r5176 (rst, clk, in, r5176_out);
	reg32 r5177 (rst, clk, in, r5177_out);
	reg32 r5178 (rst, clk, in, r5178_out);
	reg32 r5179 (rst, clk, in, r5179_out);
	reg32 r5180 (rst, clk, in, r5180_out);
	reg32 r5181 (rst, clk, in, r5181_out);
	reg32 r5182 (rst, clk, in, r5182_out);
	reg32 r5183 (rst, clk, in, r5183_out);
	reg32 r5184 (rst, clk, in, r5184_out);
	reg32 r5185 (rst, clk, in, r5185_out);
	reg32 r5186 (rst, clk, in, r5186_out);
	reg32 r5187 (rst, clk, in, r5187_out);
	reg32 r5188 (rst, clk, in, r5188_out);
	reg32 r5189 (rst, clk, in, r5189_out);
	reg32 r5190 (rst, clk, in, r5190_out);
	reg32 r5191 (rst, clk, in, r5191_out);
	reg32 r5192 (rst, clk, in, r5192_out);
	reg32 r5193 (rst, clk, in, r5193_out);
	reg32 r5194 (rst, clk, in, r5194_out);
	reg32 r5195 (rst, clk, in, r5195_out);
	reg32 r5196 (rst, clk, in, r5196_out);
	reg32 r5197 (rst, clk, in, r5197_out);
	reg32 r5198 (rst, clk, in, r5198_out);
	reg32 r5199 (rst, clk, in, r5199_out);
	reg32 r5200 (rst, clk, in, r5200_out);
	reg32 r5201 (rst, clk, in, r5201_out);
	reg32 r5202 (rst, clk, in, r5202_out);
	reg32 r5203 (rst, clk, in, r5203_out);
	reg32 r5204 (rst, clk, in, r5204_out);
	reg32 r5205 (rst, clk, in, r5205_out);
	reg32 r5206 (rst, clk, in, r5206_out);
	reg32 r5207 (rst, clk, in, r5207_out);
	reg32 r5208 (rst, clk, in, r5208_out);
	reg32 r5209 (rst, clk, in, r5209_out);
	reg32 r5210 (rst, clk, in, r5210_out);
	reg32 r5211 (rst, clk, in, r5211_out);
	reg32 r5212 (rst, clk, in, r5212_out);
	reg32 r5213 (rst, clk, in, r5213_out);
	reg32 r5214 (rst, clk, in, r5214_out);
	reg32 r5215 (rst, clk, in, r5215_out);
	reg32 r5216 (rst, clk, in, r5216_out);
	reg32 r5217 (rst, clk, in, r5217_out);
	reg32 r5218 (rst, clk, in, r5218_out);
	reg32 r5219 (rst, clk, in, r5219_out);
	reg32 r5220 (rst, clk, in, r5220_out);
	reg32 r5221 (rst, clk, in, r5221_out);
	reg32 r5222 (rst, clk, in, r5222_out);
	reg32 r5223 (rst, clk, in, r5223_out);
	reg32 r5224 (rst, clk, in, r5224_out);
	reg32 r5225 (rst, clk, in, r5225_out);
	reg32 r5226 (rst, clk, in, r5226_out);
	reg32 r5227 (rst, clk, in, r5227_out);
	reg32 r5228 (rst, clk, in, r5228_out);
	reg32 r5229 (rst, clk, in, r5229_out);
	reg32 r5230 (rst, clk, in, r5230_out);
	reg32 r5231 (rst, clk, in, r5231_out);
	reg32 r5232 (rst, clk, in, r5232_out);
	reg32 r5233 (rst, clk, in, r5233_out);
	reg32 r5234 (rst, clk, in, r5234_out);
	reg32 r5235 (rst, clk, in, r5235_out);
	reg32 r5236 (rst, clk, in, r5236_out);
	reg32 r5237 (rst, clk, in, r5237_out);
	reg32 r5238 (rst, clk, in, r5238_out);
	reg32 r5239 (rst, clk, in, r5239_out);
	reg32 r5240 (rst, clk, in, r5240_out);
	reg32 r5241 (rst, clk, in, r5241_out);
	reg32 r5242 (rst, clk, in, r5242_out);
	reg32 r5243 (rst, clk, in, r5243_out);
	reg32 r5244 (rst, clk, in, r5244_out);
	reg32 r5245 (rst, clk, in, r5245_out);
	reg32 r5246 (rst, clk, in, r5246_out);
	reg32 r5247 (rst, clk, in, r5247_out);
	reg32 r5248 (rst, clk, in, r5248_out);
	reg32 r5249 (rst, clk, in, r5249_out);
	reg32 r5250 (rst, clk, in, r5250_out);
	reg32 r5251 (rst, clk, in, r5251_out);
	reg32 r5252 (rst, clk, in, r5252_out);
	reg32 r5253 (rst, clk, in, r5253_out);
	reg32 r5254 (rst, clk, in, r5254_out);
	reg32 r5255 (rst, clk, in, r5255_out);
	reg32 r5256 (rst, clk, in, r5256_out);
	reg32 r5257 (rst, clk, in, r5257_out);
	reg32 r5258 (rst, clk, in, r5258_out);
	reg32 r5259 (rst, clk, in, r5259_out);
	reg32 r5260 (rst, clk, in, r5260_out);
	reg32 r5261 (rst, clk, in, r5261_out);
	reg32 r5262 (rst, clk, in, r5262_out);
	reg32 r5263 (rst, clk, in, r5263_out);
	reg32 r5264 (rst, clk, in, r5264_out);
	reg32 r5265 (rst, clk, in, r5265_out);
	reg32 r5266 (rst, clk, in, r5266_out);
	reg32 r5267 (rst, clk, in, r5267_out);
	reg32 r5268 (rst, clk, in, r5268_out);
	reg32 r5269 (rst, clk, in, r5269_out);
	reg32 r5270 (rst, clk, in, r5270_out);
	reg32 r5271 (rst, clk, in, r5271_out);
	reg32 r5272 (rst, clk, in, r5272_out);
	reg32 r5273 (rst, clk, in, r5273_out);
	reg32 r5274 (rst, clk, in, r5274_out);
	reg32 r5275 (rst, clk, in, r5275_out);
	reg32 r5276 (rst, clk, in, r5276_out);
	reg32 r5277 (rst, clk, in, r5277_out);
	reg32 r5278 (rst, clk, in, r5278_out);
	reg32 r5279 (rst, clk, in, r5279_out);
	reg32 r5280 (rst, clk, in, r5280_out);
	reg32 r5281 (rst, clk, in, r5281_out);
	reg32 r5282 (rst, clk, in, r5282_out);
	reg32 r5283 (rst, clk, in, r5283_out);
	reg32 r5284 (rst, clk, in, r5284_out);
	reg32 r5285 (rst, clk, in, r5285_out);
	reg32 r5286 (rst, clk, in, r5286_out);
	reg32 r5287 (rst, clk, in, r5287_out);
	reg32 r5288 (rst, clk, in, r5288_out);
	reg32 r5289 (rst, clk, in, r5289_out);
	reg32 r5290 (rst, clk, in, r5290_out);
	reg32 r5291 (rst, clk, in, r5291_out);
	reg32 r5292 (rst, clk, in, r5292_out);
	reg32 r5293 (rst, clk, in, r5293_out);
	reg32 r5294 (rst, clk, in, r5294_out);
	reg32 r5295 (rst, clk, in, r5295_out);
	reg32 r5296 (rst, clk, in, r5296_out);
	reg32 r5297 (rst, clk, in, r5297_out);
	reg32 r5298 (rst, clk, in, r5298_out);
	reg32 r5299 (rst, clk, in, r5299_out);
	reg32 r5300 (rst, clk, in, r5300_out);
	reg32 r5301 (rst, clk, in, r5301_out);
	reg32 r5302 (rst, clk, in, r5302_out);
	reg32 r5303 (rst, clk, in, r5303_out);
	reg32 r5304 (rst, clk, in, r5304_out);
	reg32 r5305 (rst, clk, in, r5305_out);
	reg32 r5306 (rst, clk, in, r5306_out);
	reg32 r5307 (rst, clk, in, r5307_out);
	reg32 r5308 (rst, clk, in, r5308_out);
	reg32 r5309 (rst, clk, in, r5309_out);
	reg32 r5310 (rst, clk, in, r5310_out);
	reg32 r5311 (rst, clk, in, r5311_out);
	reg32 r5312 (rst, clk, in, r5312_out);
	reg32 r5313 (rst, clk, in, r5313_out);
	reg32 r5314 (rst, clk, in, r5314_out);
	reg32 r5315 (rst, clk, in, r5315_out);
	reg32 r5316 (rst, clk, in, r5316_out);
	reg32 r5317 (rst, clk, in, r5317_out);
	reg32 r5318 (rst, clk, in, r5318_out);
	reg32 r5319 (rst, clk, in, r5319_out);
	reg32 r5320 (rst, clk, in, r5320_out);
	reg32 r5321 (rst, clk, in, r5321_out);
	reg32 r5322 (rst, clk, in, r5322_out);
	reg32 r5323 (rst, clk, in, r5323_out);
	reg32 r5324 (rst, clk, in, r5324_out);
	reg32 r5325 (rst, clk, in, r5325_out);
	reg32 r5326 (rst, clk, in, r5326_out);
	reg32 r5327 (rst, clk, in, r5327_out);
	reg32 r5328 (rst, clk, in, r5328_out);
	reg32 r5329 (rst, clk, in, r5329_out);
	reg32 r5330 (rst, clk, in, r5330_out);
	reg32 r5331 (rst, clk, in, r5331_out);
	reg32 r5332 (rst, clk, in, r5332_out);
	reg32 r5333 (rst, clk, in, r5333_out);
	reg32 r5334 (rst, clk, in, r5334_out);
	reg32 r5335 (rst, clk, in, r5335_out);
	reg32 r5336 (rst, clk, in, r5336_out);
	reg32 r5337 (rst, clk, in, r5337_out);
	reg32 r5338 (rst, clk, in, r5338_out);
	reg32 r5339 (rst, clk, in, r5339_out);
	reg32 r5340 (rst, clk, in, r5340_out);
	reg32 r5341 (rst, clk, in, r5341_out);
	reg32 r5342 (rst, clk, in, r5342_out);
	reg32 r5343 (rst, clk, in, r5343_out);
	reg32 r5344 (rst, clk, in, r5344_out);
	reg32 r5345 (rst, clk, in, r5345_out);
	reg32 r5346 (rst, clk, in, r5346_out);
	reg32 r5347 (rst, clk, in, r5347_out);
	reg32 r5348 (rst, clk, in, r5348_out);
	reg32 r5349 (rst, clk, in, r5349_out);
	reg32 r5350 (rst, clk, in, r5350_out);
	reg32 r5351 (rst, clk, in, r5351_out);
	reg32 r5352 (rst, clk, in, r5352_out);
	reg32 r5353 (rst, clk, in, r5353_out);
	reg32 r5354 (rst, clk, in, r5354_out);
	reg32 r5355 (rst, clk, in, r5355_out);
	reg32 r5356 (rst, clk, in, r5356_out);
	reg32 r5357 (rst, clk, in, r5357_out);
	reg32 r5358 (rst, clk, in, r5358_out);
	reg32 r5359 (rst, clk, in, r5359_out);
	reg32 r5360 (rst, clk, in, r5360_out);
	reg32 r5361 (rst, clk, in, r5361_out);
	reg32 r5362 (rst, clk, in, r5362_out);
	reg32 r5363 (rst, clk, in, r5363_out);
	reg32 r5364 (rst, clk, in, r5364_out);
	reg32 r5365 (rst, clk, in, r5365_out);
	reg32 r5366 (rst, clk, in, r5366_out);
	reg32 r5367 (rst, clk, in, r5367_out);
	reg32 r5368 (rst, clk, in, r5368_out);
	reg32 r5369 (rst, clk, in, r5369_out);
	reg32 r5370 (rst, clk, in, r5370_out);
	reg32 r5371 (rst, clk, in, r5371_out);
	reg32 r5372 (rst, clk, in, r5372_out);
	reg32 r5373 (rst, clk, in, r5373_out);
	reg32 r5374 (rst, clk, in, r5374_out);
	reg32 r5375 (rst, clk, in, r5375_out);
	reg32 r5376 (rst, clk, in, r5376_out);
	reg32 r5377 (rst, clk, in, r5377_out);
	reg32 r5378 (rst, clk, in, r5378_out);
	reg32 r5379 (rst, clk, in, r5379_out);
	reg32 r5380 (rst, clk, in, r5380_out);
	reg32 r5381 (rst, clk, in, r5381_out);
	reg32 r5382 (rst, clk, in, r5382_out);
	reg32 r5383 (rst, clk, in, r5383_out);
	reg32 r5384 (rst, clk, in, r5384_out);
	reg32 r5385 (rst, clk, in, r5385_out);
	reg32 r5386 (rst, clk, in, r5386_out);
	reg32 r5387 (rst, clk, in, r5387_out);
	reg32 r5388 (rst, clk, in, r5388_out);
	reg32 r5389 (rst, clk, in, r5389_out);
	reg32 r5390 (rst, clk, in, r5390_out);
	reg32 r5391 (rst, clk, in, r5391_out);
	reg32 r5392 (rst, clk, in, r5392_out);
	reg32 r5393 (rst, clk, in, r5393_out);
	reg32 r5394 (rst, clk, in, r5394_out);
	reg32 r5395 (rst, clk, in, r5395_out);
	reg32 r5396 (rst, clk, in, r5396_out);
	reg32 r5397 (rst, clk, in, r5397_out);
	reg32 r5398 (rst, clk, in, r5398_out);
	reg32 r5399 (rst, clk, in, r5399_out);
	reg32 r5400 (rst, clk, in, r5400_out);
	reg32 r5401 (rst, clk, in, r5401_out);
	reg32 r5402 (rst, clk, in, r5402_out);
	reg32 r5403 (rst, clk, in, r5403_out);
	reg32 r5404 (rst, clk, in, r5404_out);
	reg32 r5405 (rst, clk, in, r5405_out);
	reg32 r5406 (rst, clk, in, r5406_out);
	reg32 r5407 (rst, clk, in, r5407_out);
	reg32 r5408 (rst, clk, in, r5408_out);
	reg32 r5409 (rst, clk, in, r5409_out);
	reg32 r5410 (rst, clk, in, r5410_out);
	reg32 r5411 (rst, clk, in, r5411_out);
	reg32 r5412 (rst, clk, in, r5412_out);
	reg32 r5413 (rst, clk, in, r5413_out);
	reg32 r5414 (rst, clk, in, r5414_out);
	reg32 r5415 (rst, clk, in, r5415_out);
	reg32 r5416 (rst, clk, in, r5416_out);
	reg32 r5417 (rst, clk, in, r5417_out);
	reg32 r5418 (rst, clk, in, r5418_out);
	reg32 r5419 (rst, clk, in, r5419_out);
	reg32 r5420 (rst, clk, in, r5420_out);
	reg32 r5421 (rst, clk, in, r5421_out);
	reg32 r5422 (rst, clk, in, r5422_out);
	reg32 r5423 (rst, clk, in, r5423_out);
	reg32 r5424 (rst, clk, in, r5424_out);
	reg32 r5425 (rst, clk, in, r5425_out);
	reg32 r5426 (rst, clk, in, r5426_out);
	reg32 r5427 (rst, clk, in, r5427_out);
	reg32 r5428 (rst, clk, in, r5428_out);
	reg32 r5429 (rst, clk, in, r5429_out);
	reg32 r5430 (rst, clk, in, r5430_out);
	reg32 r5431 (rst, clk, in, r5431_out);
	reg32 r5432 (rst, clk, in, r5432_out);
	reg32 r5433 (rst, clk, in, r5433_out);
	reg32 r5434 (rst, clk, in, r5434_out);
	reg32 r5435 (rst, clk, in, r5435_out);
	reg32 r5436 (rst, clk, in, r5436_out);
	reg32 r5437 (rst, clk, in, r5437_out);
	reg32 r5438 (rst, clk, in, r5438_out);
	reg32 r5439 (rst, clk, in, r5439_out);
	reg32 r5440 (rst, clk, in, r5440_out);
	reg32 r5441 (rst, clk, in, r5441_out);
	reg32 r5442 (rst, clk, in, r5442_out);
	reg32 r5443 (rst, clk, in, r5443_out);
	reg32 r5444 (rst, clk, in, r5444_out);
	reg32 r5445 (rst, clk, in, r5445_out);
	reg32 r5446 (rst, clk, in, r5446_out);
	reg32 r5447 (rst, clk, in, r5447_out);
	reg32 r5448 (rst, clk, in, r5448_out);
	reg32 r5449 (rst, clk, in, r5449_out);
	reg32 r5450 (rst, clk, in, r5450_out);
	reg32 r5451 (rst, clk, in, r5451_out);
	reg32 r5452 (rst, clk, in, r5452_out);
	reg32 r5453 (rst, clk, in, r5453_out);
	reg32 r5454 (rst, clk, in, r5454_out);
	reg32 r5455 (rst, clk, in, r5455_out);
	reg32 r5456 (rst, clk, in, r5456_out);
	reg32 r5457 (rst, clk, in, r5457_out);
	reg32 r5458 (rst, clk, in, r5458_out);
	reg32 r5459 (rst, clk, in, r5459_out);
	reg32 r5460 (rst, clk, in, r5460_out);
	reg32 r5461 (rst, clk, in, r5461_out);
	reg32 r5462 (rst, clk, in, r5462_out);
	reg32 r5463 (rst, clk, in, r5463_out);
	reg32 r5464 (rst, clk, in, r5464_out);
	reg32 r5465 (rst, clk, in, r5465_out);
	reg32 r5466 (rst, clk, in, r5466_out);
	reg32 r5467 (rst, clk, in, r5467_out);
	reg32 r5468 (rst, clk, in, r5468_out);
	reg32 r5469 (rst, clk, in, r5469_out);
	reg32 r5470 (rst, clk, in, r5470_out);
	reg32 r5471 (rst, clk, in, r5471_out);
	reg32 r5472 (rst, clk, in, r5472_out);
	reg32 r5473 (rst, clk, in, r5473_out);
	reg32 r5474 (rst, clk, in, r5474_out);
	reg32 r5475 (rst, clk, in, r5475_out);
	reg32 r5476 (rst, clk, in, r5476_out);
	reg32 r5477 (rst, clk, in, r5477_out);
	reg32 r5478 (rst, clk, in, r5478_out);
	reg32 r5479 (rst, clk, in, r5479_out);
	reg32 r5480 (rst, clk, in, r5480_out);
	reg32 r5481 (rst, clk, in, r5481_out);
	reg32 r5482 (rst, clk, in, r5482_out);
	reg32 r5483 (rst, clk, in, r5483_out);
	reg32 r5484 (rst, clk, in, r5484_out);
	reg32 r5485 (rst, clk, in, r5485_out);
	reg32 r5486 (rst, clk, in, r5486_out);
	reg32 r5487 (rst, clk, in, r5487_out);
	reg32 r5488 (rst, clk, in, r5488_out);
	reg32 r5489 (rst, clk, in, r5489_out);
	reg32 r5490 (rst, clk, in, r5490_out);
	reg32 r5491 (rst, clk, in, r5491_out);
	reg32 r5492 (rst, clk, in, r5492_out);
	reg32 r5493 (rst, clk, in, r5493_out);
	reg32 r5494 (rst, clk, in, r5494_out);
	reg32 r5495 (rst, clk, in, r5495_out);
	reg32 r5496 (rst, clk, in, r5496_out);
	reg32 r5497 (rst, clk, in, r5497_out);
	reg32 r5498 (rst, clk, in, r5498_out);
	reg32 r5499 (rst, clk, in, r5499_out);
	reg32 r5500 (rst, clk, in, r5500_out);
	reg32 r5501 (rst, clk, in, r5501_out);
	reg32 r5502 (rst, clk, in, r5502_out);
	reg32 r5503 (rst, clk, in, r5503_out);
	reg32 r5504 (rst, clk, in, r5504_out);
	reg32 r5505 (rst, clk, in, r5505_out);
	reg32 r5506 (rst, clk, in, r5506_out);
	reg32 r5507 (rst, clk, in, r5507_out);
	reg32 r5508 (rst, clk, in, r5508_out);
	reg32 r5509 (rst, clk, in, r5509_out);
	reg32 r5510 (rst, clk, in, r5510_out);
	reg32 r5511 (rst, clk, in, r5511_out);
	reg32 r5512 (rst, clk, in, r5512_out);
	reg32 r5513 (rst, clk, in, r5513_out);
	reg32 r5514 (rst, clk, in, r5514_out);
	reg32 r5515 (rst, clk, in, r5515_out);
	reg32 r5516 (rst, clk, in, r5516_out);
	reg32 r5517 (rst, clk, in, r5517_out);
	reg32 r5518 (rst, clk, in, r5518_out);
	reg32 r5519 (rst, clk, in, r5519_out);
	reg32 r5520 (rst, clk, in, r5520_out);
	reg32 r5521 (rst, clk, in, r5521_out);
	reg32 r5522 (rst, clk, in, r5522_out);
	reg32 r5523 (rst, clk, in, r5523_out);
	reg32 r5524 (rst, clk, in, r5524_out);
	reg32 r5525 (rst, clk, in, r5525_out);
	reg32 r5526 (rst, clk, in, r5526_out);
	reg32 r5527 (rst, clk, in, r5527_out);
	reg32 r5528 (rst, clk, in, r5528_out);
	reg32 r5529 (rst, clk, in, r5529_out);
	reg32 r5530 (rst, clk, in, r5530_out);
	reg32 r5531 (rst, clk, in, r5531_out);
	reg32 r5532 (rst, clk, in, r5532_out);
	reg32 r5533 (rst, clk, in, r5533_out);
	reg32 r5534 (rst, clk, in, r5534_out);
	reg32 r5535 (rst, clk, in, r5535_out);
	reg32 r5536 (rst, clk, in, r5536_out);
	reg32 r5537 (rst, clk, in, r5537_out);
	reg32 r5538 (rst, clk, in, r5538_out);
	reg32 r5539 (rst, clk, in, r5539_out);
	reg32 r5540 (rst, clk, in, r5540_out);
	reg32 r5541 (rst, clk, in, r5541_out);
	reg32 r5542 (rst, clk, in, r5542_out);
	reg32 r5543 (rst, clk, in, r5543_out);
	reg32 r5544 (rst, clk, in, r5544_out);
	reg32 r5545 (rst, clk, in, r5545_out);
	reg32 r5546 (rst, clk, in, r5546_out);
	reg32 r5547 (rst, clk, in, r5547_out);
	reg32 r5548 (rst, clk, in, r5548_out);
	reg32 r5549 (rst, clk, in, r5549_out);
	reg32 r5550 (rst, clk, in, r5550_out);
	reg32 r5551 (rst, clk, in, r5551_out);
	reg32 r5552 (rst, clk, in, r5552_out);
	reg32 r5553 (rst, clk, in, r5553_out);
	reg32 r5554 (rst, clk, in, r5554_out);
	reg32 r5555 (rst, clk, in, r5555_out);
	reg32 r5556 (rst, clk, in, r5556_out);
	reg32 r5557 (rst, clk, in, r5557_out);
	reg32 r5558 (rst, clk, in, r5558_out);
	reg32 r5559 (rst, clk, in, r5559_out);
	reg32 r5560 (rst, clk, in, r5560_out);
	reg32 r5561 (rst, clk, in, r5561_out);
	reg32 r5562 (rst, clk, in, r5562_out);
	reg32 r5563 (rst, clk, in, r5563_out);
	reg32 r5564 (rst, clk, in, r5564_out);
	reg32 r5565 (rst, clk, in, r5565_out);
	reg32 r5566 (rst, clk, in, r5566_out);
	reg32 r5567 (rst, clk, in, r5567_out);
	reg32 r5568 (rst, clk, in, r5568_out);
	reg32 r5569 (rst, clk, in, r5569_out);
	reg32 r5570 (rst, clk, in, r5570_out);
	reg32 r5571 (rst, clk, in, r5571_out);
	reg32 r5572 (rst, clk, in, r5572_out);
	reg32 r5573 (rst, clk, in, r5573_out);
	reg32 r5574 (rst, clk, in, r5574_out);
	reg32 r5575 (rst, clk, in, r5575_out);
	reg32 r5576 (rst, clk, in, r5576_out);
	reg32 r5577 (rst, clk, in, r5577_out);
	reg32 r5578 (rst, clk, in, r5578_out);
	reg32 r5579 (rst, clk, in, r5579_out);
	reg32 r5580 (rst, clk, in, r5580_out);
	reg32 r5581 (rst, clk, in, r5581_out);
	reg32 r5582 (rst, clk, in, r5582_out);
	reg32 r5583 (rst, clk, in, r5583_out);
	reg32 r5584 (rst, clk, in, r5584_out);
	reg32 r5585 (rst, clk, in, r5585_out);
	reg32 r5586 (rst, clk, in, r5586_out);
	reg32 r5587 (rst, clk, in, r5587_out);
	reg32 r5588 (rst, clk, in, r5588_out);
	reg32 r5589 (rst, clk, in, r5589_out);
	reg32 r5590 (rst, clk, in, r5590_out);
	reg32 r5591 (rst, clk, in, r5591_out);
	reg32 r5592 (rst, clk, in, r5592_out);
	reg32 r5593 (rst, clk, in, r5593_out);
	reg32 r5594 (rst, clk, in, r5594_out);
	reg32 r5595 (rst, clk, in, r5595_out);
	reg32 r5596 (rst, clk, in, r5596_out);
	reg32 r5597 (rst, clk, in, r5597_out);
	reg32 r5598 (rst, clk, in, r5598_out);
	reg32 r5599 (rst, clk, in, r5599_out);
	reg32 r5600 (rst, clk, in, r5600_out);
	reg32 r5601 (rst, clk, in, r5601_out);
	reg32 r5602 (rst, clk, in, r5602_out);
	reg32 r5603 (rst, clk, in, r5603_out);
	reg32 r5604 (rst, clk, in, r5604_out);
	reg32 r5605 (rst, clk, in, r5605_out);
	reg32 r5606 (rst, clk, in, r5606_out);
	reg32 r5607 (rst, clk, in, r5607_out);
	reg32 r5608 (rst, clk, in, r5608_out);
	reg32 r5609 (rst, clk, in, r5609_out);
	reg32 r5610 (rst, clk, in, r5610_out);
	reg32 r5611 (rst, clk, in, r5611_out);
	reg32 r5612 (rst, clk, in, r5612_out);
	reg32 r5613 (rst, clk, in, r5613_out);
	reg32 r5614 (rst, clk, in, r5614_out);
	reg32 r5615 (rst, clk, in, r5615_out);
	reg32 r5616 (rst, clk, in, r5616_out);
	reg32 r5617 (rst, clk, in, r5617_out);
	reg32 r5618 (rst, clk, in, r5618_out);
	reg32 r5619 (rst, clk, in, r5619_out);
	reg32 r5620 (rst, clk, in, r5620_out);
	reg32 r5621 (rst, clk, in, r5621_out);
	reg32 r5622 (rst, clk, in, r5622_out);
	reg32 r5623 (rst, clk, in, r5623_out);
	reg32 r5624 (rst, clk, in, r5624_out);
	reg32 r5625 (rst, clk, in, r5625_out);
	reg32 r5626 (rst, clk, in, r5626_out);
	reg32 r5627 (rst, clk, in, r5627_out);
	reg32 r5628 (rst, clk, in, r5628_out);
	reg32 r5629 (rst, clk, in, r5629_out);
	reg32 r5630 (rst, clk, in, r5630_out);
	reg32 r5631 (rst, clk, in, r5631_out);
	reg32 r5632 (rst, clk, in, r5632_out);
	reg32 r5633 (rst, clk, in, r5633_out);
	reg32 r5634 (rst, clk, in, r5634_out);
	reg32 r5635 (rst, clk, in, r5635_out);
	reg32 r5636 (rst, clk, in, r5636_out);
	reg32 r5637 (rst, clk, in, r5637_out);
	reg32 r5638 (rst, clk, in, r5638_out);
	reg32 r5639 (rst, clk, in, r5639_out);
	reg32 r5640 (rst, clk, in, r5640_out);
	reg32 r5641 (rst, clk, in, r5641_out);
	reg32 r5642 (rst, clk, in, r5642_out);
	reg32 r5643 (rst, clk, in, r5643_out);
	reg32 r5644 (rst, clk, in, r5644_out);
	reg32 r5645 (rst, clk, in, r5645_out);
	reg32 r5646 (rst, clk, in, r5646_out);
	reg32 r5647 (rst, clk, in, r5647_out);
	reg32 r5648 (rst, clk, in, r5648_out);
	reg32 r5649 (rst, clk, in, r5649_out);
	reg32 r5650 (rst, clk, in, r5650_out);
	reg32 r5651 (rst, clk, in, r5651_out);
	reg32 r5652 (rst, clk, in, r5652_out);
	reg32 r5653 (rst, clk, in, r5653_out);
	reg32 r5654 (rst, clk, in, r5654_out);
	reg32 r5655 (rst, clk, in, r5655_out);
	reg32 r5656 (rst, clk, in, r5656_out);
	reg32 r5657 (rst, clk, in, r5657_out);
	reg32 r5658 (rst, clk, in, r5658_out);
	reg32 r5659 (rst, clk, in, r5659_out);
	reg32 r5660 (rst, clk, in, r5660_out);
	reg32 r5661 (rst, clk, in, r5661_out);
	reg32 r5662 (rst, clk, in, r5662_out);
	reg32 r5663 (rst, clk, in, r5663_out);
	reg32 r5664 (rst, clk, in, r5664_out);
	reg32 r5665 (rst, clk, in, r5665_out);
	reg32 r5666 (rst, clk, in, r5666_out);
	reg32 r5667 (rst, clk, in, r5667_out);
	reg32 r5668 (rst, clk, in, r5668_out);
	reg32 r5669 (rst, clk, in, r5669_out);
	reg32 r5670 (rst, clk, in, r5670_out);
	reg32 r5671 (rst, clk, in, r5671_out);
	reg32 r5672 (rst, clk, in, r5672_out);
	reg32 r5673 (rst, clk, in, r5673_out);
	reg32 r5674 (rst, clk, in, r5674_out);
	reg32 r5675 (rst, clk, in, r5675_out);
	reg32 r5676 (rst, clk, in, r5676_out);
	reg32 r5677 (rst, clk, in, r5677_out);
	reg32 r5678 (rst, clk, in, r5678_out);
	reg32 r5679 (rst, clk, in, r5679_out);
	reg32 r5680 (rst, clk, in, r5680_out);
	reg32 r5681 (rst, clk, in, r5681_out);
	reg32 r5682 (rst, clk, in, r5682_out);
	reg32 r5683 (rst, clk, in, r5683_out);
	reg32 r5684 (rst, clk, in, r5684_out);
	reg32 r5685 (rst, clk, in, r5685_out);
	reg32 r5686 (rst, clk, in, r5686_out);
	reg32 r5687 (rst, clk, in, r5687_out);
	reg32 r5688 (rst, clk, in, r5688_out);
	reg32 r5689 (rst, clk, in, r5689_out);
	reg32 r5690 (rst, clk, in, r5690_out);
	reg32 r5691 (rst, clk, in, r5691_out);
	reg32 r5692 (rst, clk, in, r5692_out);
	reg32 r5693 (rst, clk, in, r5693_out);
	reg32 r5694 (rst, clk, in, r5694_out);
	reg32 r5695 (rst, clk, in, r5695_out);
	reg32 r5696 (rst, clk, in, r5696_out);
	reg32 r5697 (rst, clk, in, r5697_out);
	reg32 r5698 (rst, clk, in, r5698_out);
	reg32 r5699 (rst, clk, in, r5699_out);
	reg32 r5700 (rst, clk, in, r5700_out);
	reg32 r5701 (rst, clk, in, r5701_out);
	reg32 r5702 (rst, clk, in, r5702_out);
	reg32 r5703 (rst, clk, in, r5703_out);
	reg32 r5704 (rst, clk, in, r5704_out);
	reg32 r5705 (rst, clk, in, r5705_out);
	reg32 r5706 (rst, clk, in, r5706_out);
	reg32 r5707 (rst, clk, in, r5707_out);
	reg32 r5708 (rst, clk, in, r5708_out);
	reg32 r5709 (rst, clk, in, r5709_out);
	reg32 r5710 (rst, clk, in, r5710_out);
	reg32 r5711 (rst, clk, in, r5711_out);
	reg32 r5712 (rst, clk, in, r5712_out);
	reg32 r5713 (rst, clk, in, r5713_out);
	reg32 r5714 (rst, clk, in, r5714_out);
	reg32 r5715 (rst, clk, in, r5715_out);
	reg32 r5716 (rst, clk, in, r5716_out);
	reg32 r5717 (rst, clk, in, r5717_out);
	reg32 r5718 (rst, clk, in, r5718_out);
	reg32 r5719 (rst, clk, in, r5719_out);
	reg32 r5720 (rst, clk, in, r5720_out);
	reg32 r5721 (rst, clk, in, r5721_out);
	reg32 r5722 (rst, clk, in, r5722_out);
	reg32 r5723 (rst, clk, in, r5723_out);
	reg32 r5724 (rst, clk, in, r5724_out);
	reg32 r5725 (rst, clk, in, r5725_out);
	reg32 r5726 (rst, clk, in, r5726_out);
	reg32 r5727 (rst, clk, in, r5727_out);
	reg32 r5728 (rst, clk, in, r5728_out);
	reg32 r5729 (rst, clk, in, r5729_out);
	reg32 r5730 (rst, clk, in, r5730_out);
	reg32 r5731 (rst, clk, in, r5731_out);
	reg32 r5732 (rst, clk, in, r5732_out);
	reg32 r5733 (rst, clk, in, r5733_out);
	reg32 r5734 (rst, clk, in, r5734_out);
	reg32 r5735 (rst, clk, in, r5735_out);
	reg32 r5736 (rst, clk, in, r5736_out);
	reg32 r5737 (rst, clk, in, r5737_out);
	reg32 r5738 (rst, clk, in, r5738_out);
	reg32 r5739 (rst, clk, in, r5739_out);
	reg32 r5740 (rst, clk, in, r5740_out);
	reg32 r5741 (rst, clk, in, r5741_out);
	reg32 r5742 (rst, clk, in, r5742_out);
	reg32 r5743 (rst, clk, in, r5743_out);
	reg32 r5744 (rst, clk, in, r5744_out);
	reg32 r5745 (rst, clk, in, r5745_out);
	reg32 r5746 (rst, clk, in, r5746_out);
	reg32 r5747 (rst, clk, in, r5747_out);
	reg32 r5748 (rst, clk, in, r5748_out);
	reg32 r5749 (rst, clk, in, r5749_out);
	reg32 r5750 (rst, clk, in, r5750_out);
	reg32 r5751 (rst, clk, in, r5751_out);
	reg32 r5752 (rst, clk, in, r5752_out);
	reg32 r5753 (rst, clk, in, r5753_out);
	reg32 r5754 (rst, clk, in, r5754_out);
	reg32 r5755 (rst, clk, in, r5755_out);
	reg32 r5756 (rst, clk, in, r5756_out);
	reg32 r5757 (rst, clk, in, r5757_out);
	reg32 r5758 (rst, clk, in, r5758_out);
	reg32 r5759 (rst, clk, in, r5759_out);
	reg32 r5760 (rst, clk, in, r5760_out);
	reg32 r5761 (rst, clk, in, r5761_out);
	reg32 r5762 (rst, clk, in, r5762_out);
	reg32 r5763 (rst, clk, in, r5763_out);
	reg32 r5764 (rst, clk, in, r5764_out);
	reg32 r5765 (rst, clk, in, r5765_out);
	reg32 r5766 (rst, clk, in, r5766_out);
	reg32 r5767 (rst, clk, in, r5767_out);
	reg32 r5768 (rst, clk, in, r5768_out);
	reg32 r5769 (rst, clk, in, r5769_out);
	reg32 r5770 (rst, clk, in, r5770_out);
	reg32 r5771 (rst, clk, in, r5771_out);
	reg32 r5772 (rst, clk, in, r5772_out);
	reg32 r5773 (rst, clk, in, r5773_out);
	reg32 r5774 (rst, clk, in, r5774_out);
	reg32 r5775 (rst, clk, in, r5775_out);
	reg32 r5776 (rst, clk, in, r5776_out);
	reg32 r5777 (rst, clk, in, r5777_out);
	reg32 r5778 (rst, clk, in, r5778_out);
	reg32 r5779 (rst, clk, in, r5779_out);
	reg32 r5780 (rst, clk, in, r5780_out);
	reg32 r5781 (rst, clk, in, r5781_out);
	reg32 r5782 (rst, clk, in, r5782_out);
	reg32 r5783 (rst, clk, in, r5783_out);
	reg32 r5784 (rst, clk, in, r5784_out);
	reg32 r5785 (rst, clk, in, r5785_out);
	reg32 r5786 (rst, clk, in, r5786_out);
	reg32 r5787 (rst, clk, in, r5787_out);
	reg32 r5788 (rst, clk, in, r5788_out);
	reg32 r5789 (rst, clk, in, r5789_out);
	reg32 r5790 (rst, clk, in, r5790_out);
	reg32 r5791 (rst, clk, in, r5791_out);
	reg32 r5792 (rst, clk, in, r5792_out);
	reg32 r5793 (rst, clk, in, r5793_out);
	reg32 r5794 (rst, clk, in, r5794_out);
	reg32 r5795 (rst, clk, in, r5795_out);
	reg32 r5796 (rst, clk, in, r5796_out);
	reg32 r5797 (rst, clk, in, r5797_out);
	reg32 r5798 (rst, clk, in, r5798_out);
	reg32 r5799 (rst, clk, in, r5799_out);
	reg32 r5800 (rst, clk, in, r5800_out);
	reg32 r5801 (rst, clk, in, r5801_out);
	reg32 r5802 (rst, clk, in, r5802_out);
	reg32 r5803 (rst, clk, in, r5803_out);
	reg32 r5804 (rst, clk, in, r5804_out);
	reg32 r5805 (rst, clk, in, r5805_out);
	reg32 r5806 (rst, clk, in, r5806_out);
	reg32 r5807 (rst, clk, in, r5807_out);
	reg32 r5808 (rst, clk, in, r5808_out);
	reg32 r5809 (rst, clk, in, r5809_out);
	reg32 r5810 (rst, clk, in, r5810_out);
	reg32 r5811 (rst, clk, in, r5811_out);
	reg32 r5812 (rst, clk, in, r5812_out);
	reg32 r5813 (rst, clk, in, r5813_out);
	reg32 r5814 (rst, clk, in, r5814_out);
	reg32 r5815 (rst, clk, in, r5815_out);
	reg32 r5816 (rst, clk, in, r5816_out);
	reg32 r5817 (rst, clk, in, r5817_out);
	reg32 r5818 (rst, clk, in, r5818_out);
	reg32 r5819 (rst, clk, in, r5819_out);
	reg32 r5820 (rst, clk, in, r5820_out);
	reg32 r5821 (rst, clk, in, r5821_out);
	reg32 r5822 (rst, clk, in, r5822_out);
	reg32 r5823 (rst, clk, in, r5823_out);
	reg32 r5824 (rst, clk, in, r5824_out);
	reg32 r5825 (rst, clk, in, r5825_out);
	reg32 r5826 (rst, clk, in, r5826_out);
	reg32 r5827 (rst, clk, in, r5827_out);
	reg32 r5828 (rst, clk, in, r5828_out);
	reg32 r5829 (rst, clk, in, r5829_out);
	reg32 r5830 (rst, clk, in, r5830_out);
	reg32 r5831 (rst, clk, in, r5831_out);
	reg32 r5832 (rst, clk, in, r5832_out);
	reg32 r5833 (rst, clk, in, r5833_out);
	reg32 r5834 (rst, clk, in, r5834_out);
	reg32 r5835 (rst, clk, in, r5835_out);
	reg32 r5836 (rst, clk, in, r5836_out);
	reg32 r5837 (rst, clk, in, r5837_out);
	reg32 r5838 (rst, clk, in, r5838_out);
	reg32 r5839 (rst, clk, in, r5839_out);
	reg32 r5840 (rst, clk, in, r5840_out);
	reg32 r5841 (rst, clk, in, r5841_out);
	reg32 r5842 (rst, clk, in, r5842_out);
	reg32 r5843 (rst, clk, in, r5843_out);
	reg32 r5844 (rst, clk, in, r5844_out);
	reg32 r5845 (rst, clk, in, r5845_out);
	reg32 r5846 (rst, clk, in, r5846_out);
	reg32 r5847 (rst, clk, in, r5847_out);
	reg32 r5848 (rst, clk, in, r5848_out);
	reg32 r5849 (rst, clk, in, r5849_out);
	reg32 r5850 (rst, clk, in, r5850_out);
	reg32 r5851 (rst, clk, in, r5851_out);
	reg32 r5852 (rst, clk, in, r5852_out);
	reg32 r5853 (rst, clk, in, r5853_out);
	reg32 r5854 (rst, clk, in, r5854_out);
	reg32 r5855 (rst, clk, in, r5855_out);
	reg32 r5856 (rst, clk, in, r5856_out);
	reg32 r5857 (rst, clk, in, r5857_out);
	reg32 r5858 (rst, clk, in, r5858_out);
	reg32 r5859 (rst, clk, in, r5859_out);
	reg32 r5860 (rst, clk, in, r5860_out);
	reg32 r5861 (rst, clk, in, r5861_out);
	reg32 r5862 (rst, clk, in, r5862_out);
	reg32 r5863 (rst, clk, in, r5863_out);
	reg32 r5864 (rst, clk, in, r5864_out);
	reg32 r5865 (rst, clk, in, r5865_out);
	reg32 r5866 (rst, clk, in, r5866_out);
	reg32 r5867 (rst, clk, in, r5867_out);
	reg32 r5868 (rst, clk, in, r5868_out);
	reg32 r5869 (rst, clk, in, r5869_out);
	reg32 r5870 (rst, clk, in, r5870_out);
	reg32 r5871 (rst, clk, in, r5871_out);
	reg32 r5872 (rst, clk, in, r5872_out);
	reg32 r5873 (rst, clk, in, r5873_out);
	reg32 r5874 (rst, clk, in, r5874_out);
	reg32 r5875 (rst, clk, in, r5875_out);
	reg32 r5876 (rst, clk, in, r5876_out);
	reg32 r5877 (rst, clk, in, r5877_out);
	reg32 r5878 (rst, clk, in, r5878_out);
	reg32 r5879 (rst, clk, in, r5879_out);
	reg32 r5880 (rst, clk, in, r5880_out);
	reg32 r5881 (rst, clk, in, r5881_out);
	reg32 r5882 (rst, clk, in, r5882_out);
	reg32 r5883 (rst, clk, in, r5883_out);
	reg32 r5884 (rst, clk, in, r5884_out);
	reg32 r5885 (rst, clk, in, r5885_out);
	reg32 r5886 (rst, clk, in, r5886_out);
	reg32 r5887 (rst, clk, in, r5887_out);
	reg32 r5888 (rst, clk, in, r5888_out);
	reg32 r5889 (rst, clk, in, r5889_out);
	reg32 r5890 (rst, clk, in, r5890_out);
	reg32 r5891 (rst, clk, in, r5891_out);
	reg32 r5892 (rst, clk, in, r5892_out);
	reg32 r5893 (rst, clk, in, r5893_out);
	reg32 r5894 (rst, clk, in, r5894_out);
	reg32 r5895 (rst, clk, in, r5895_out);
	reg32 r5896 (rst, clk, in, r5896_out);
	reg32 r5897 (rst, clk, in, r5897_out);
	reg32 r5898 (rst, clk, in, r5898_out);
	reg32 r5899 (rst, clk, in, r5899_out);
	reg32 r5900 (rst, clk, in, r5900_out);
	reg32 r5901 (rst, clk, in, r5901_out);
	reg32 r5902 (rst, clk, in, r5902_out);
	reg32 r5903 (rst, clk, in, r5903_out);
	reg32 r5904 (rst, clk, in, r5904_out);
	reg32 r5905 (rst, clk, in, r5905_out);
	reg32 r5906 (rst, clk, in, r5906_out);
	reg32 r5907 (rst, clk, in, r5907_out);
	reg32 r5908 (rst, clk, in, r5908_out);
	reg32 r5909 (rst, clk, in, r5909_out);
	reg32 r5910 (rst, clk, in, r5910_out);
	reg32 r5911 (rst, clk, in, r5911_out);
	reg32 r5912 (rst, clk, in, r5912_out);
	reg32 r5913 (rst, clk, in, r5913_out);
	reg32 r5914 (rst, clk, in, r5914_out);
	reg32 r5915 (rst, clk, in, r5915_out);
	reg32 r5916 (rst, clk, in, r5916_out);
	reg32 r5917 (rst, clk, in, r5917_out);
	reg32 r5918 (rst, clk, in, r5918_out);
	reg32 r5919 (rst, clk, in, r5919_out);
	reg32 r5920 (rst, clk, in, r5920_out);
	reg32 r5921 (rst, clk, in, r5921_out);
	reg32 r5922 (rst, clk, in, r5922_out);
	reg32 r5923 (rst, clk, in, r5923_out);
	reg32 r5924 (rst, clk, in, r5924_out);
	reg32 r5925 (rst, clk, in, r5925_out);
	reg32 r5926 (rst, clk, in, r5926_out);
	reg32 r5927 (rst, clk, in, r5927_out);
	reg32 r5928 (rst, clk, in, r5928_out);
	reg32 r5929 (rst, clk, in, r5929_out);
	reg32 r5930 (rst, clk, in, r5930_out);
	reg32 r5931 (rst, clk, in, r5931_out);
	reg32 r5932 (rst, clk, in, r5932_out);
	reg32 r5933 (rst, clk, in, r5933_out);
	reg32 r5934 (rst, clk, in, r5934_out);
	reg32 r5935 (rst, clk, in, r5935_out);
	reg32 r5936 (rst, clk, in, r5936_out);
	reg32 r5937 (rst, clk, in, r5937_out);
	reg32 r5938 (rst, clk, in, r5938_out);
	reg32 r5939 (rst, clk, in, r5939_out);
	reg32 r5940 (rst, clk, in, r5940_out);
	reg32 r5941 (rst, clk, in, r5941_out);
	reg32 r5942 (rst, clk, in, r5942_out);
	reg32 r5943 (rst, clk, in, r5943_out);
	reg32 r5944 (rst, clk, in, r5944_out);
	reg32 r5945 (rst, clk, in, r5945_out);
	reg32 r5946 (rst, clk, in, r5946_out);
	reg32 r5947 (rst, clk, in, r5947_out);
	reg32 r5948 (rst, clk, in, r5948_out);
	reg32 r5949 (rst, clk, in, r5949_out);
	reg32 r5950 (rst, clk, in, r5950_out);
	reg32 r5951 (rst, clk, in, r5951_out);
	reg32 r5952 (rst, clk, in, r5952_out);
	reg32 r5953 (rst, clk, in, r5953_out);
	reg32 r5954 (rst, clk, in, r5954_out);
	reg32 r5955 (rst, clk, in, r5955_out);
	reg32 r5956 (rst, clk, in, r5956_out);
	reg32 r5957 (rst, clk, in, r5957_out);
	reg32 r5958 (rst, clk, in, r5958_out);
	reg32 r5959 (rst, clk, in, r5959_out);
	reg32 r5960 (rst, clk, in, r5960_out);
	reg32 r5961 (rst, clk, in, r5961_out);
	reg32 r5962 (rst, clk, in, r5962_out);
	reg32 r5963 (rst, clk, in, r5963_out);
	reg32 r5964 (rst, clk, in, r5964_out);
	reg32 r5965 (rst, clk, in, r5965_out);
	reg32 r5966 (rst, clk, in, r5966_out);
	reg32 r5967 (rst, clk, in, r5967_out);
	reg32 r5968 (rst, clk, in, r5968_out);
	reg32 r5969 (rst, clk, in, r5969_out);
	reg32 r5970 (rst, clk, in, r5970_out);
	reg32 r5971 (rst, clk, in, r5971_out);
	reg32 r5972 (rst, clk, in, r5972_out);
	reg32 r5973 (rst, clk, in, r5973_out);
	reg32 r5974 (rst, clk, in, r5974_out);
	reg32 r5975 (rst, clk, in, r5975_out);
	reg32 r5976 (rst, clk, in, r5976_out);
	reg32 r5977 (rst, clk, in, r5977_out);
	reg32 r5978 (rst, clk, in, r5978_out);
	reg32 r5979 (rst, clk, in, r5979_out);
	reg32 r5980 (rst, clk, in, r5980_out);
	reg32 r5981 (rst, clk, in, r5981_out);
	reg32 r5982 (rst, clk, in, r5982_out);
	reg32 r5983 (rst, clk, in, r5983_out);
	reg32 r5984 (rst, clk, in, r5984_out);
	reg32 r5985 (rst, clk, in, r5985_out);
	reg32 r5986 (rst, clk, in, r5986_out);
	reg32 r5987 (rst, clk, in, r5987_out);
	reg32 r5988 (rst, clk, in, r5988_out);
	reg32 r5989 (rst, clk, in, r5989_out);
	reg32 r5990 (rst, clk, in, r5990_out);
	reg32 r5991 (rst, clk, in, r5991_out);
	reg32 r5992 (rst, clk, in, r5992_out);
	reg32 r5993 (rst, clk, in, r5993_out);
	reg32 r5994 (rst, clk, in, r5994_out);
	reg32 r5995 (rst, clk, in, r5995_out);
	reg32 r5996 (rst, clk, in, r5996_out);
	reg32 r5997 (rst, clk, in, r5997_out);
	reg32 r5998 (rst, clk, in, r5998_out);
	reg32 r5999 (rst, clk, in, r5999_out);
	reg32 r6000 (rst, clk, in, r6000_out);
	reg32 r6001 (rst, clk, in, r6001_out);
	reg32 r6002 (rst, clk, in, r6002_out);
	reg32 r6003 (rst, clk, in, r6003_out);
	reg32 r6004 (rst, clk, in, r6004_out);
	reg32 r6005 (rst, clk, in, r6005_out);
	reg32 r6006 (rst, clk, in, r6006_out);
	reg32 r6007 (rst, clk, in, r6007_out);
	reg32 r6008 (rst, clk, in, r6008_out);
	reg32 r6009 (rst, clk, in, r6009_out);
	reg32 r6010 (rst, clk, in, r6010_out);
	reg32 r6011 (rst, clk, in, r6011_out);
	reg32 r6012 (rst, clk, in, r6012_out);
	reg32 r6013 (rst, clk, in, r6013_out);
	reg32 r6014 (rst, clk, in, r6014_out);
	reg32 r6015 (rst, clk, in, r6015_out);
	reg32 r6016 (rst, clk, in, r6016_out);
	reg32 r6017 (rst, clk, in, r6017_out);
	reg32 r6018 (rst, clk, in, r6018_out);
	reg32 r6019 (rst, clk, in, r6019_out);
	reg32 r6020 (rst, clk, in, r6020_out);
	reg32 r6021 (rst, clk, in, r6021_out);
	reg32 r6022 (rst, clk, in, r6022_out);
	reg32 r6023 (rst, clk, in, r6023_out);
	reg32 r6024 (rst, clk, in, r6024_out);
	reg32 r6025 (rst, clk, in, r6025_out);
	reg32 r6026 (rst, clk, in, r6026_out);
	reg32 r6027 (rst, clk, in, r6027_out);
	reg32 r6028 (rst, clk, in, r6028_out);
	reg32 r6029 (rst, clk, in, r6029_out);
	reg32 r6030 (rst, clk, in, r6030_out);
	reg32 r6031 (rst, clk, in, r6031_out);
	reg32 r6032 (rst, clk, in, r6032_out);
	reg32 r6033 (rst, clk, in, r6033_out);
	reg32 r6034 (rst, clk, in, r6034_out);
	reg32 r6035 (rst, clk, in, r6035_out);
	reg32 r6036 (rst, clk, in, r6036_out);
	reg32 r6037 (rst, clk, in, r6037_out);
	reg32 r6038 (rst, clk, in, r6038_out);
	reg32 r6039 (rst, clk, in, r6039_out);
	reg32 r6040 (rst, clk, in, r6040_out);
	reg32 r6041 (rst, clk, in, r6041_out);
	reg32 r6042 (rst, clk, in, r6042_out);
	reg32 r6043 (rst, clk, in, r6043_out);
	reg32 r6044 (rst, clk, in, r6044_out);
	reg32 r6045 (rst, clk, in, r6045_out);
	reg32 r6046 (rst, clk, in, r6046_out);
	reg32 r6047 (rst, clk, in, r6047_out);
	reg32 r6048 (rst, clk, in, r6048_out);
	reg32 r6049 (rst, clk, in, r6049_out);
	reg32 r6050 (rst, clk, in, r6050_out);
	reg32 r6051 (rst, clk, in, r6051_out);
	reg32 r6052 (rst, clk, in, r6052_out);
	reg32 r6053 (rst, clk, in, r6053_out);
	reg32 r6054 (rst, clk, in, r6054_out);
	reg32 r6055 (rst, clk, in, r6055_out);
	reg32 r6056 (rst, clk, in, r6056_out);
	reg32 r6057 (rst, clk, in, r6057_out);
	reg32 r6058 (rst, clk, in, r6058_out);
	reg32 r6059 (rst, clk, in, r6059_out);
	reg32 r6060 (rst, clk, in, r6060_out);
	reg32 r6061 (rst, clk, in, r6061_out);
	reg32 r6062 (rst, clk, in, r6062_out);
	reg32 r6063 (rst, clk, in, r6063_out);
	reg32 r6064 (rst, clk, in, r6064_out);
	reg32 r6065 (rst, clk, in, r6065_out);
	reg32 r6066 (rst, clk, in, r6066_out);
	reg32 r6067 (rst, clk, in, r6067_out);
	reg32 r6068 (rst, clk, in, r6068_out);
	reg32 r6069 (rst, clk, in, r6069_out);
	reg32 r6070 (rst, clk, in, r6070_out);
	reg32 r6071 (rst, clk, in, r6071_out);
	reg32 r6072 (rst, clk, in, r6072_out);
	reg32 r6073 (rst, clk, in, r6073_out);
	reg32 r6074 (rst, clk, in, r6074_out);
	reg32 r6075 (rst, clk, in, r6075_out);
	reg32 r6076 (rst, clk, in, r6076_out);
	reg32 r6077 (rst, clk, in, r6077_out);
	reg32 r6078 (rst, clk, in, r6078_out);
	reg32 r6079 (rst, clk, in, r6079_out);
	reg32 r6080 (rst, clk, in, r6080_out);
	reg32 r6081 (rst, clk, in, r6081_out);
	reg32 r6082 (rst, clk, in, r6082_out);
	reg32 r6083 (rst, clk, in, r6083_out);
	reg32 r6084 (rst, clk, in, r6084_out);
	reg32 r6085 (rst, clk, in, r6085_out);
	reg32 r6086 (rst, clk, in, r6086_out);
	reg32 r6087 (rst, clk, in, r6087_out);
	reg32 r6088 (rst, clk, in, r6088_out);
	reg32 r6089 (rst, clk, in, r6089_out);
	reg32 r6090 (rst, clk, in, r6090_out);
	reg32 r6091 (rst, clk, in, r6091_out);
	reg32 r6092 (rst, clk, in, r6092_out);
	reg32 r6093 (rst, clk, in, r6093_out);
	reg32 r6094 (rst, clk, in, r6094_out);
	reg32 r6095 (rst, clk, in, r6095_out);
	reg32 r6096 (rst, clk, in, r6096_out);
	reg32 r6097 (rst, clk, in, r6097_out);
	reg32 r6098 (rst, clk, in, r6098_out);
	reg32 r6099 (rst, clk, in, r6099_out);
	reg32 r6100 (rst, clk, in, r6100_out);
	reg32 r6101 (rst, clk, in, r6101_out);
	reg32 r6102 (rst, clk, in, r6102_out);
	reg32 r6103 (rst, clk, in, r6103_out);
	reg32 r6104 (rst, clk, in, r6104_out);
	reg32 r6105 (rst, clk, in, r6105_out);
	reg32 r6106 (rst, clk, in, r6106_out);
	reg32 r6107 (rst, clk, in, r6107_out);
	reg32 r6108 (rst, clk, in, r6108_out);
	reg32 r6109 (rst, clk, in, r6109_out);
	reg32 r6110 (rst, clk, in, r6110_out);
	reg32 r6111 (rst, clk, in, r6111_out);
	reg32 r6112 (rst, clk, in, r6112_out);
	reg32 r6113 (rst, clk, in, r6113_out);
	reg32 r6114 (rst, clk, in, r6114_out);
	reg32 r6115 (rst, clk, in, r6115_out);
	reg32 r6116 (rst, clk, in, r6116_out);
	reg32 r6117 (rst, clk, in, r6117_out);
	reg32 r6118 (rst, clk, in, r6118_out);
	reg32 r6119 (rst, clk, in, r6119_out);
	reg32 r6120 (rst, clk, in, r6120_out);
	reg32 r6121 (rst, clk, in, r6121_out);
	reg32 r6122 (rst, clk, in, r6122_out);
	reg32 r6123 (rst, clk, in, r6123_out);
	reg32 r6124 (rst, clk, in, r6124_out);
	reg32 r6125 (rst, clk, in, r6125_out);
	reg32 r6126 (rst, clk, in, r6126_out);
	reg32 r6127 (rst, clk, in, r6127_out);
	reg32 r6128 (rst, clk, in, r6128_out);
	reg32 r6129 (rst, clk, in, r6129_out);
	reg32 r6130 (rst, clk, in, r6130_out);
	reg32 r6131 (rst, clk, in, r6131_out);
	reg32 r6132 (rst, clk, in, r6132_out);
	reg32 r6133 (rst, clk, in, r6133_out);
	reg32 r6134 (rst, clk, in, r6134_out);
	reg32 r6135 (rst, clk, in, r6135_out);
	reg32 r6136 (rst, clk, in, r6136_out);
	reg32 r6137 (rst, clk, in, r6137_out);
	reg32 r6138 (rst, clk, in, r6138_out);
	reg32 r6139 (rst, clk, in, r6139_out);
	reg32 r6140 (rst, clk, in, r6140_out);
	reg32 r6141 (rst, clk, in, r6141_out);
	reg32 r6142 (rst, clk, in, r6142_out);
	reg32 r6143 (rst, clk, in, r6143_out);
	reg32 r6144 (rst, clk, in, r6144_out);
	reg32 r6145 (rst, clk, in, r6145_out);
	reg32 r6146 (rst, clk, in, r6146_out);
	reg32 r6147 (rst, clk, in, r6147_out);
	reg32 r6148 (rst, clk, in, r6148_out);
	reg32 r6149 (rst, clk, in, r6149_out);
	reg32 r6150 (rst, clk, in, r6150_out);
	reg32 r6151 (rst, clk, in, r6151_out);
	reg32 r6152 (rst, clk, in, r6152_out);
	reg32 r6153 (rst, clk, in, r6153_out);
	reg32 r6154 (rst, clk, in, r6154_out);
	reg32 r6155 (rst, clk, in, r6155_out);
	reg32 r6156 (rst, clk, in, r6156_out);
	reg32 r6157 (rst, clk, in, r6157_out);
	reg32 r6158 (rst, clk, in, r6158_out);
	reg32 r6159 (rst, clk, in, r6159_out);
	reg32 r6160 (rst, clk, in, r6160_out);
	reg32 r6161 (rst, clk, in, r6161_out);
	reg32 r6162 (rst, clk, in, r6162_out);
	reg32 r6163 (rst, clk, in, r6163_out);
	reg32 r6164 (rst, clk, in, r6164_out);
	reg32 r6165 (rst, clk, in, r6165_out);
	reg32 r6166 (rst, clk, in, r6166_out);
	reg32 r6167 (rst, clk, in, r6167_out);
	reg32 r6168 (rst, clk, in, r6168_out);
	reg32 r6169 (rst, clk, in, r6169_out);
	reg32 r6170 (rst, clk, in, r6170_out);
	reg32 r6171 (rst, clk, in, r6171_out);
	reg32 r6172 (rst, clk, in, r6172_out);
	reg32 r6173 (rst, clk, in, r6173_out);
	reg32 r6174 (rst, clk, in, r6174_out);
	reg32 r6175 (rst, clk, in, r6175_out);
	reg32 r6176 (rst, clk, in, r6176_out);
	reg32 r6177 (rst, clk, in, r6177_out);
	reg32 r6178 (rst, clk, in, r6178_out);
	reg32 r6179 (rst, clk, in, r6179_out);
	reg32 r6180 (rst, clk, in, r6180_out);
	reg32 r6181 (rst, clk, in, r6181_out);
	reg32 r6182 (rst, clk, in, r6182_out);
	reg32 r6183 (rst, clk, in, r6183_out);
	reg32 r6184 (rst, clk, in, r6184_out);
	reg32 r6185 (rst, clk, in, r6185_out);
	reg32 r6186 (rst, clk, in, r6186_out);
	reg32 r6187 (rst, clk, in, r6187_out);
	reg32 r6188 (rst, clk, in, r6188_out);
	reg32 r6189 (rst, clk, in, r6189_out);
	reg32 r6190 (rst, clk, in, r6190_out);
	reg32 r6191 (rst, clk, in, r6191_out);
	reg32 r6192 (rst, clk, in, r6192_out);
	reg32 r6193 (rst, clk, in, r6193_out);
	reg32 r6194 (rst, clk, in, r6194_out);
	reg32 r6195 (rst, clk, in, r6195_out);
	reg32 r6196 (rst, clk, in, r6196_out);
	reg32 r6197 (rst, clk, in, r6197_out);
	reg32 r6198 (rst, clk, in, r6198_out);
	reg32 r6199 (rst, clk, in, r6199_out);
	reg32 r6200 (rst, clk, in, r6200_out);
	reg32 r6201 (rst, clk, in, r6201_out);
	reg32 r6202 (rst, clk, in, r6202_out);
	reg32 r6203 (rst, clk, in, r6203_out);
	reg32 r6204 (rst, clk, in, r6204_out);
	reg32 r6205 (rst, clk, in, r6205_out);
	reg32 r6206 (rst, clk, in, r6206_out);
	reg32 r6207 (rst, clk, in, r6207_out);
	reg32 r6208 (rst, clk, in, r6208_out);
	reg32 r6209 (rst, clk, in, r6209_out);
	reg32 r6210 (rst, clk, in, r6210_out);
	reg32 r6211 (rst, clk, in, r6211_out);
	reg32 r6212 (rst, clk, in, r6212_out);
	reg32 r6213 (rst, clk, in, r6213_out);
	reg32 r6214 (rst, clk, in, r6214_out);
	reg32 r6215 (rst, clk, in, r6215_out);
	reg32 r6216 (rst, clk, in, r6216_out);
	reg32 r6217 (rst, clk, in, r6217_out);
	reg32 r6218 (rst, clk, in, r6218_out);
	reg32 r6219 (rst, clk, in, r6219_out);
	reg32 r6220 (rst, clk, in, r6220_out);
	reg32 r6221 (rst, clk, in, r6221_out);
	reg32 r6222 (rst, clk, in, r6222_out);
	reg32 r6223 (rst, clk, in, r6223_out);
	reg32 r6224 (rst, clk, in, r6224_out);
	reg32 r6225 (rst, clk, in, r6225_out);
	reg32 r6226 (rst, clk, in, r6226_out);
	reg32 r6227 (rst, clk, in, r6227_out);
	reg32 r6228 (rst, clk, in, r6228_out);
	reg32 r6229 (rst, clk, in, r6229_out);
	reg32 r6230 (rst, clk, in, r6230_out);
	reg32 r6231 (rst, clk, in, r6231_out);
	reg32 r6232 (rst, clk, in, r6232_out);
	reg32 r6233 (rst, clk, in, r6233_out);
	reg32 r6234 (rst, clk, in, r6234_out);
	reg32 r6235 (rst, clk, in, r6235_out);
	reg32 r6236 (rst, clk, in, r6236_out);
	reg32 r6237 (rst, clk, in, r6237_out);
	reg32 r6238 (rst, clk, in, r6238_out);
	reg32 r6239 (rst, clk, in, r6239_out);
	reg32 r6240 (rst, clk, in, r6240_out);
	reg32 r6241 (rst, clk, in, r6241_out);
	reg32 r6242 (rst, clk, in, r6242_out);
	reg32 r6243 (rst, clk, in, r6243_out);
	reg32 r6244 (rst, clk, in, r6244_out);
	reg32 r6245 (rst, clk, in, r6245_out);
	reg32 r6246 (rst, clk, in, r6246_out);
	reg32 r6247 (rst, clk, in, r6247_out);
	reg32 r6248 (rst, clk, in, r6248_out);
	reg32 r6249 (rst, clk, in, r6249_out);
	reg32 r6250 (rst, clk, in, r6250_out);
	reg32 r6251 (rst, clk, in, r6251_out);
	reg32 r6252 (rst, clk, in, r6252_out);
	reg32 r6253 (rst, clk, in, r6253_out);
	reg32 r6254 (rst, clk, in, r6254_out);
	reg32 r6255 (rst, clk, in, r6255_out);
	reg32 r6256 (rst, clk, in, r6256_out);
	reg32 r6257 (rst, clk, in, r6257_out);
	reg32 r6258 (rst, clk, in, r6258_out);
	reg32 r6259 (rst, clk, in, r6259_out);
	reg32 r6260 (rst, clk, in, r6260_out);
	reg32 r6261 (rst, clk, in, r6261_out);
	reg32 r6262 (rst, clk, in, r6262_out);
	reg32 r6263 (rst, clk, in, r6263_out);
	reg32 r6264 (rst, clk, in, r6264_out);
	reg32 r6265 (rst, clk, in, r6265_out);
	reg32 r6266 (rst, clk, in, r6266_out);
	reg32 r6267 (rst, clk, in, r6267_out);
	reg32 r6268 (rst, clk, in, r6268_out);
	reg32 r6269 (rst, clk, in, r6269_out);
	reg32 r6270 (rst, clk, in, r6270_out);
	reg32 r6271 (rst, clk, in, r6271_out);
	reg32 r6272 (rst, clk, in, r6272_out);
	reg32 r6273 (rst, clk, in, r6273_out);
	reg32 r6274 (rst, clk, in, r6274_out);
	reg32 r6275 (rst, clk, in, r6275_out);
	reg32 r6276 (rst, clk, in, r6276_out);
	reg32 r6277 (rst, clk, in, r6277_out);
	reg32 r6278 (rst, clk, in, r6278_out);
	reg32 r6279 (rst, clk, in, r6279_out);
	reg32 r6280 (rst, clk, in, r6280_out);
	reg32 r6281 (rst, clk, in, r6281_out);
	reg32 r6282 (rst, clk, in, r6282_out);
	reg32 r6283 (rst, clk, in, r6283_out);
	reg32 r6284 (rst, clk, in, r6284_out);
	reg32 r6285 (rst, clk, in, r6285_out);
	reg32 r6286 (rst, clk, in, r6286_out);
	reg32 r6287 (rst, clk, in, r6287_out);
	reg32 r6288 (rst, clk, in, r6288_out);
	reg32 r6289 (rst, clk, in, r6289_out);
	reg32 r6290 (rst, clk, in, r6290_out);
	reg32 r6291 (rst, clk, in, r6291_out);
	reg32 r6292 (rst, clk, in, r6292_out);
	reg32 r6293 (rst, clk, in, r6293_out);
	reg32 r6294 (rst, clk, in, r6294_out);
	reg32 r6295 (rst, clk, in, r6295_out);
	reg32 r6296 (rst, clk, in, r6296_out);
	reg32 r6297 (rst, clk, in, r6297_out);
	reg32 r6298 (rst, clk, in, r6298_out);
	reg32 r6299 (rst, clk, in, r6299_out);
	reg32 r6300 (rst, clk, in, r6300_out);
	reg32 r6301 (rst, clk, in, r6301_out);
	reg32 r6302 (rst, clk, in, r6302_out);
	reg32 r6303 (rst, clk, in, r6303_out);
	reg32 r6304 (rst, clk, in, r6304_out);
	reg32 r6305 (rst, clk, in, r6305_out);
	reg32 r6306 (rst, clk, in, r6306_out);
	reg32 r6307 (rst, clk, in, r6307_out);
	reg32 r6308 (rst, clk, in, r6308_out);
	reg32 r6309 (rst, clk, in, r6309_out);
	reg32 r6310 (rst, clk, in, r6310_out);
	reg32 r6311 (rst, clk, in, r6311_out);
	reg32 r6312 (rst, clk, in, r6312_out);
	reg32 r6313 (rst, clk, in, r6313_out);
	reg32 r6314 (rst, clk, in, r6314_out);
	reg32 r6315 (rst, clk, in, r6315_out);
	reg32 r6316 (rst, clk, in, r6316_out);
	reg32 r6317 (rst, clk, in, r6317_out);
	reg32 r6318 (rst, clk, in, r6318_out);
	reg32 r6319 (rst, clk, in, r6319_out);
	reg32 r6320 (rst, clk, in, r6320_out);
	reg32 r6321 (rst, clk, in, r6321_out);
	reg32 r6322 (rst, clk, in, r6322_out);
	reg32 r6323 (rst, clk, in, r6323_out);
	reg32 r6324 (rst, clk, in, r6324_out);
	reg32 r6325 (rst, clk, in, r6325_out);
	reg32 r6326 (rst, clk, in, r6326_out);
	reg32 r6327 (rst, clk, in, r6327_out);
	reg32 r6328 (rst, clk, in, r6328_out);
	reg32 r6329 (rst, clk, in, r6329_out);
	reg32 r6330 (rst, clk, in, r6330_out);
	reg32 r6331 (rst, clk, in, r6331_out);
	reg32 r6332 (rst, clk, in, r6332_out);
	reg32 r6333 (rst, clk, in, r6333_out);
	reg32 r6334 (rst, clk, in, r6334_out);
	reg32 r6335 (rst, clk, in, r6335_out);
	reg32 r6336 (rst, clk, in, r6336_out);
	reg32 r6337 (rst, clk, in, r6337_out);
	reg32 r6338 (rst, clk, in, r6338_out);
	reg32 r6339 (rst, clk, in, r6339_out);
	reg32 r6340 (rst, clk, in, r6340_out);
	reg32 r6341 (rst, clk, in, r6341_out);
	reg32 r6342 (rst, clk, in, r6342_out);
	reg32 r6343 (rst, clk, in, r6343_out);
	reg32 r6344 (rst, clk, in, r6344_out);
	reg32 r6345 (rst, clk, in, r6345_out);
	reg32 r6346 (rst, clk, in, r6346_out);
	reg32 r6347 (rst, clk, in, r6347_out);
	reg32 r6348 (rst, clk, in, r6348_out);
	reg32 r6349 (rst, clk, in, r6349_out);
	reg32 r6350 (rst, clk, in, r6350_out);
	reg32 r6351 (rst, clk, in, r6351_out);
	reg32 r6352 (rst, clk, in, r6352_out);
	reg32 r6353 (rst, clk, in, r6353_out);
	reg32 r6354 (rst, clk, in, r6354_out);
	reg32 r6355 (rst, clk, in, r6355_out);
	reg32 r6356 (rst, clk, in, r6356_out);
	reg32 r6357 (rst, clk, in, r6357_out);
	reg32 r6358 (rst, clk, in, r6358_out);
	reg32 r6359 (rst, clk, in, r6359_out);
	reg32 r6360 (rst, clk, in, r6360_out);
	reg32 r6361 (rst, clk, in, r6361_out);
	reg32 r6362 (rst, clk, in, r6362_out);
	reg32 r6363 (rst, clk, in, r6363_out);
	reg32 r6364 (rst, clk, in, r6364_out);
	reg32 r6365 (rst, clk, in, r6365_out);
	reg32 r6366 (rst, clk, in, r6366_out);
	reg32 r6367 (rst, clk, in, r6367_out);
	reg32 r6368 (rst, clk, in, r6368_out);
	reg32 r6369 (rst, clk, in, r6369_out);
	reg32 r6370 (rst, clk, in, r6370_out);
	reg32 r6371 (rst, clk, in, r6371_out);
	reg32 r6372 (rst, clk, in, r6372_out);
	reg32 r6373 (rst, clk, in, r6373_out);
	reg32 r6374 (rst, clk, in, r6374_out);
	reg32 r6375 (rst, clk, in, r6375_out);
	reg32 r6376 (rst, clk, in, r6376_out);
	reg32 r6377 (rst, clk, in, r6377_out);
	reg32 r6378 (rst, clk, in, r6378_out);
	reg32 r6379 (rst, clk, in, r6379_out);
	reg32 r6380 (rst, clk, in, r6380_out);
	reg32 r6381 (rst, clk, in, r6381_out);
	reg32 r6382 (rst, clk, in, r6382_out);
	reg32 r6383 (rst, clk, in, r6383_out);
	reg32 r6384 (rst, clk, in, r6384_out);
	reg32 r6385 (rst, clk, in, r6385_out);
	reg32 r6386 (rst, clk, in, r6386_out);
	reg32 r6387 (rst, clk, in, r6387_out);
	reg32 r6388 (rst, clk, in, r6388_out);
	reg32 r6389 (rst, clk, in, r6389_out);
	reg32 r6390 (rst, clk, in, r6390_out);
	reg32 r6391 (rst, clk, in, r6391_out);
	reg32 r6392 (rst, clk, in, r6392_out);
	reg32 r6393 (rst, clk, in, r6393_out);
	reg32 r6394 (rst, clk, in, r6394_out);
	reg32 r6395 (rst, clk, in, r6395_out);
	reg32 r6396 (rst, clk, in, r6396_out);
	reg32 r6397 (rst, clk, in, r6397_out);
	reg32 r6398 (rst, clk, in, r6398_out);
	reg32 r6399 (rst, clk, in, r6399_out);
	reg32 r6400 (rst, clk, in, r6400_out);
	reg32 r6401 (rst, clk, in, r6401_out);
	reg32 r6402 (rst, clk, in, r6402_out);
	reg32 r6403 (rst, clk, in, r6403_out);
	reg32 r6404 (rst, clk, in, r6404_out);
	reg32 r6405 (rst, clk, in, r6405_out);
	reg32 r6406 (rst, clk, in, r6406_out);
	reg32 r6407 (rst, clk, in, r6407_out);
	reg32 r6408 (rst, clk, in, r6408_out);
	reg32 r6409 (rst, clk, in, r6409_out);
	reg32 r6410 (rst, clk, in, r6410_out);
	reg32 r6411 (rst, clk, in, r6411_out);
	reg32 r6412 (rst, clk, in, r6412_out);
	reg32 r6413 (rst, clk, in, r6413_out);
	reg32 r6414 (rst, clk, in, r6414_out);
	reg32 r6415 (rst, clk, in, r6415_out);
	reg32 r6416 (rst, clk, in, r6416_out);
	reg32 r6417 (rst, clk, in, r6417_out);
	reg32 r6418 (rst, clk, in, r6418_out);
	reg32 r6419 (rst, clk, in, r6419_out);
	reg32 r6420 (rst, clk, in, r6420_out);
	reg32 r6421 (rst, clk, in, r6421_out);
	reg32 r6422 (rst, clk, in, r6422_out);
	reg32 r6423 (rst, clk, in, r6423_out);
	reg32 r6424 (rst, clk, in, r6424_out);
	reg32 r6425 (rst, clk, in, r6425_out);
	reg32 r6426 (rst, clk, in, r6426_out);
	reg32 r6427 (rst, clk, in, r6427_out);
	reg32 r6428 (rst, clk, in, r6428_out);
	reg32 r6429 (rst, clk, in, r6429_out);
	reg32 r6430 (rst, clk, in, r6430_out);
	reg32 r6431 (rst, clk, in, r6431_out);
	reg32 r6432 (rst, clk, in, r6432_out);
	reg32 r6433 (rst, clk, in, r6433_out);
	reg32 r6434 (rst, clk, in, r6434_out);
	reg32 r6435 (rst, clk, in, r6435_out);
	reg32 r6436 (rst, clk, in, r6436_out);
	reg32 r6437 (rst, clk, in, r6437_out);
	reg32 r6438 (rst, clk, in, r6438_out);
	reg32 r6439 (rst, clk, in, r6439_out);
	reg32 r6440 (rst, clk, in, r6440_out);
	reg32 r6441 (rst, clk, in, r6441_out);
	reg32 r6442 (rst, clk, in, r6442_out);
	reg32 r6443 (rst, clk, in, r6443_out);
	reg32 r6444 (rst, clk, in, r6444_out);
	reg32 r6445 (rst, clk, in, r6445_out);
	reg32 r6446 (rst, clk, in, r6446_out);
	reg32 r6447 (rst, clk, in, r6447_out);
	reg32 r6448 (rst, clk, in, r6448_out);
	reg32 r6449 (rst, clk, in, r6449_out);
	reg32 r6450 (rst, clk, in, r6450_out);
	reg32 r6451 (rst, clk, in, r6451_out);
	reg32 r6452 (rst, clk, in, r6452_out);
	reg32 r6453 (rst, clk, in, r6453_out);
	reg32 r6454 (rst, clk, in, r6454_out);
	reg32 r6455 (rst, clk, in, r6455_out);
	reg32 r6456 (rst, clk, in, r6456_out);
	reg32 r6457 (rst, clk, in, r6457_out);
	reg32 r6458 (rst, clk, in, r6458_out);
	reg32 r6459 (rst, clk, in, r6459_out);
	reg32 r6460 (rst, clk, in, r6460_out);
	reg32 r6461 (rst, clk, in, r6461_out);
	reg32 r6462 (rst, clk, in, r6462_out);
	reg32 r6463 (rst, clk, in, r6463_out);
	reg32 r6464 (rst, clk, in, r6464_out);
	reg32 r6465 (rst, clk, in, r6465_out);
	reg32 r6466 (rst, clk, in, r6466_out);
	reg32 r6467 (rst, clk, in, r6467_out);
	reg32 r6468 (rst, clk, in, r6468_out);
	reg32 r6469 (rst, clk, in, r6469_out);
	reg32 r6470 (rst, clk, in, r6470_out);
	reg32 r6471 (rst, clk, in, r6471_out);
	reg32 r6472 (rst, clk, in, r6472_out);
	reg32 r6473 (rst, clk, in, r6473_out);
	reg32 r6474 (rst, clk, in, r6474_out);
	reg32 r6475 (rst, clk, in, r6475_out);
	reg32 r6476 (rst, clk, in, r6476_out);
	reg32 r6477 (rst, clk, in, r6477_out);
	reg32 r6478 (rst, clk, in, r6478_out);
	reg32 r6479 (rst, clk, in, r6479_out);
	reg32 r6480 (rst, clk, in, r6480_out);
	reg32 r6481 (rst, clk, in, r6481_out);
	reg32 r6482 (rst, clk, in, r6482_out);
	reg32 r6483 (rst, clk, in, r6483_out);
	reg32 r6484 (rst, clk, in, r6484_out);
	reg32 r6485 (rst, clk, in, r6485_out);
	reg32 r6486 (rst, clk, in, r6486_out);
	reg32 r6487 (rst, clk, in, r6487_out);
	reg32 r6488 (rst, clk, in, r6488_out);
	reg32 r6489 (rst, clk, in, r6489_out);
	reg32 r6490 (rst, clk, in, r6490_out);
	reg32 r6491 (rst, clk, in, r6491_out);
	reg32 r6492 (rst, clk, in, r6492_out);
	reg32 r6493 (rst, clk, in, r6493_out);
	reg32 r6494 (rst, clk, in, r6494_out);
	reg32 r6495 (rst, clk, in, r6495_out);
	reg32 r6496 (rst, clk, in, r6496_out);
	reg32 r6497 (rst, clk, in, r6497_out);
	reg32 r6498 (rst, clk, in, r6498_out);
	reg32 r6499 (rst, clk, in, r6499_out);
	reg32 r6500 (rst, clk, in, r6500_out);
	reg32 r6501 (rst, clk, in, r6501_out);
	reg32 r6502 (rst, clk, in, r6502_out);
	reg32 r6503 (rst, clk, in, r6503_out);
	reg32 r6504 (rst, clk, in, r6504_out);
	reg32 r6505 (rst, clk, in, r6505_out);
	reg32 r6506 (rst, clk, in, r6506_out);
	reg32 r6507 (rst, clk, in, r6507_out);
	reg32 r6508 (rst, clk, in, r6508_out);
	reg32 r6509 (rst, clk, in, r6509_out);
	reg32 r6510 (rst, clk, in, r6510_out);
	reg32 r6511 (rst, clk, in, r6511_out);
	reg32 r6512 (rst, clk, in, r6512_out);
	reg32 r6513 (rst, clk, in, r6513_out);
	reg32 r6514 (rst, clk, in, r6514_out);
	reg32 r6515 (rst, clk, in, r6515_out);
	reg32 r6516 (rst, clk, in, r6516_out);
	reg32 r6517 (rst, clk, in, r6517_out);
	reg32 r6518 (rst, clk, in, r6518_out);
	reg32 r6519 (rst, clk, in, r6519_out);
	reg32 r6520 (rst, clk, in, r6520_out);
	reg32 r6521 (rst, clk, in, r6521_out);
	reg32 r6522 (rst, clk, in, r6522_out);
	reg32 r6523 (rst, clk, in, r6523_out);
	reg32 r6524 (rst, clk, in, r6524_out);
	reg32 r6525 (rst, clk, in, r6525_out);
	reg32 r6526 (rst, clk, in, r6526_out);
	reg32 r6527 (rst, clk, in, r6527_out);
	reg32 r6528 (rst, clk, in, r6528_out);
	reg32 r6529 (rst, clk, in, r6529_out);
	reg32 r6530 (rst, clk, in, r6530_out);
	reg32 r6531 (rst, clk, in, r6531_out);
	reg32 r6532 (rst, clk, in, r6532_out);
	reg32 r6533 (rst, clk, in, r6533_out);
	reg32 r6534 (rst, clk, in, r6534_out);
	reg32 r6535 (rst, clk, in, r6535_out);
	reg32 r6536 (rst, clk, in, r6536_out);
	reg32 r6537 (rst, clk, in, r6537_out);
	reg32 r6538 (rst, clk, in, r6538_out);
	reg32 r6539 (rst, clk, in, r6539_out);
	reg32 r6540 (rst, clk, in, r6540_out);
	reg32 r6541 (rst, clk, in, r6541_out);
	reg32 r6542 (rst, clk, in, r6542_out);
	reg32 r6543 (rst, clk, in, r6543_out);
	reg32 r6544 (rst, clk, in, r6544_out);
	reg32 r6545 (rst, clk, in, r6545_out);
	reg32 r6546 (rst, clk, in, r6546_out);
	reg32 r6547 (rst, clk, in, r6547_out);
	reg32 r6548 (rst, clk, in, r6548_out);
	reg32 r6549 (rst, clk, in, r6549_out);
	reg32 r6550 (rst, clk, in, r6550_out);
	reg32 r6551 (rst, clk, in, r6551_out);
	reg32 r6552 (rst, clk, in, r6552_out);
	reg32 r6553 (rst, clk, in, r6553_out);
	reg32 r6554 (rst, clk, in, r6554_out);
	reg32 r6555 (rst, clk, in, r6555_out);
	reg32 r6556 (rst, clk, in, r6556_out);
	reg32 r6557 (rst, clk, in, r6557_out);
	reg32 r6558 (rst, clk, in, r6558_out);
	reg32 r6559 (rst, clk, in, r6559_out);
	reg32 r6560 (rst, clk, in, r6560_out);
	reg32 r6561 (rst, clk, in, r6561_out);
	reg32 r6562 (rst, clk, in, r6562_out);
	reg32 r6563 (rst, clk, in, r6563_out);
	reg32 r6564 (rst, clk, in, r6564_out);
	reg32 r6565 (rst, clk, in, r6565_out);
	reg32 r6566 (rst, clk, in, r6566_out);
	reg32 r6567 (rst, clk, in, r6567_out);
	reg32 r6568 (rst, clk, in, r6568_out);
	reg32 r6569 (rst, clk, in, r6569_out);
	reg32 r6570 (rst, clk, in, r6570_out);
	reg32 r6571 (rst, clk, in, r6571_out);
	reg32 r6572 (rst, clk, in, r6572_out);
	reg32 r6573 (rst, clk, in, r6573_out);
	reg32 r6574 (rst, clk, in, r6574_out);
	reg32 r6575 (rst, clk, in, r6575_out);
	reg32 r6576 (rst, clk, in, r6576_out);
	reg32 r6577 (rst, clk, in, r6577_out);
	reg32 r6578 (rst, clk, in, r6578_out);
	reg32 r6579 (rst, clk, in, r6579_out);
	reg32 r6580 (rst, clk, in, r6580_out);
	reg32 r6581 (rst, clk, in, r6581_out);
	reg32 r6582 (rst, clk, in, r6582_out);
	reg32 r6583 (rst, clk, in, r6583_out);
	reg32 r6584 (rst, clk, in, r6584_out);
	reg32 r6585 (rst, clk, in, r6585_out);
	reg32 r6586 (rst, clk, in, r6586_out);
	reg32 r6587 (rst, clk, in, r6587_out);
	reg32 r6588 (rst, clk, in, r6588_out);
	reg32 r6589 (rst, clk, in, r6589_out);
	reg32 r6590 (rst, clk, in, r6590_out);
	reg32 r6591 (rst, clk, in, r6591_out);
	reg32 r6592 (rst, clk, in, r6592_out);
	reg32 r6593 (rst, clk, in, r6593_out);
	reg32 r6594 (rst, clk, in, r6594_out);
	reg32 r6595 (rst, clk, in, r6595_out);
	reg32 r6596 (rst, clk, in, r6596_out);
	reg32 r6597 (rst, clk, in, r6597_out);
	reg32 r6598 (rst, clk, in, r6598_out);
	reg32 r6599 (rst, clk, in, r6599_out);
	reg32 r6600 (rst, clk, in, r6600_out);
	reg32 r6601 (rst, clk, in, r6601_out);
	reg32 r6602 (rst, clk, in, r6602_out);
	reg32 r6603 (rst, clk, in, r6603_out);
	reg32 r6604 (rst, clk, in, r6604_out);
	reg32 r6605 (rst, clk, in, r6605_out);
	reg32 r6606 (rst, clk, in, r6606_out);
	reg32 r6607 (rst, clk, in, r6607_out);
	reg32 r6608 (rst, clk, in, r6608_out);
	reg32 r6609 (rst, clk, in, r6609_out);
	reg32 r6610 (rst, clk, in, r6610_out);
	reg32 r6611 (rst, clk, in, r6611_out);
	reg32 r6612 (rst, clk, in, r6612_out);
	reg32 r6613 (rst, clk, in, r6613_out);
	reg32 r6614 (rst, clk, in, r6614_out);
	reg32 r6615 (rst, clk, in, r6615_out);
	reg32 r6616 (rst, clk, in, r6616_out);
	reg32 r6617 (rst, clk, in, r6617_out);
	reg32 r6618 (rst, clk, in, r6618_out);
	reg32 r6619 (rst, clk, in, r6619_out);
	reg32 r6620 (rst, clk, in, r6620_out);
	reg32 r6621 (rst, clk, in, r6621_out);
	reg32 r6622 (rst, clk, in, r6622_out);
	reg32 r6623 (rst, clk, in, r6623_out);
	reg32 r6624 (rst, clk, in, r6624_out);
	reg32 r6625 (rst, clk, in, r6625_out);
	reg32 r6626 (rst, clk, in, r6626_out);
	reg32 r6627 (rst, clk, in, r6627_out);
	reg32 r6628 (rst, clk, in, r6628_out);
	reg32 r6629 (rst, clk, in, r6629_out);
	reg32 r6630 (rst, clk, in, r6630_out);
	reg32 r6631 (rst, clk, in, r6631_out);
	reg32 r6632 (rst, clk, in, r6632_out);
	reg32 r6633 (rst, clk, in, r6633_out);
	reg32 r6634 (rst, clk, in, r6634_out);
	reg32 r6635 (rst, clk, in, r6635_out);
	reg32 r6636 (rst, clk, in, r6636_out);
	reg32 r6637 (rst, clk, in, r6637_out);
	reg32 r6638 (rst, clk, in, r6638_out);
	reg32 r6639 (rst, clk, in, r6639_out);
	reg32 r6640 (rst, clk, in, r6640_out);
	reg32 r6641 (rst, clk, in, r6641_out);
	reg32 r6642 (rst, clk, in, r6642_out);
	reg32 r6643 (rst, clk, in, r6643_out);
	reg32 r6644 (rst, clk, in, r6644_out);
	reg32 r6645 (rst, clk, in, r6645_out);
	reg32 r6646 (rst, clk, in, r6646_out);
	reg32 r6647 (rst, clk, in, r6647_out);
	reg32 r6648 (rst, clk, in, r6648_out);
	reg32 r6649 (rst, clk, in, r6649_out);
	reg32 r6650 (rst, clk, in, r6650_out);
	reg32 r6651 (rst, clk, in, r6651_out);
	reg32 r6652 (rst, clk, in, r6652_out);
	reg32 r6653 (rst, clk, in, r6653_out);
	reg32 r6654 (rst, clk, in, r6654_out);
	reg32 r6655 (rst, clk, in, r6655_out);
	reg32 r6656 (rst, clk, in, r6656_out);
	reg32 r6657 (rst, clk, in, r6657_out);
	reg32 r6658 (rst, clk, in, r6658_out);
	reg32 r6659 (rst, clk, in, r6659_out);
	reg32 r6660 (rst, clk, in, r6660_out);
	reg32 r6661 (rst, clk, in, r6661_out);
	reg32 r6662 (rst, clk, in, r6662_out);
	reg32 r6663 (rst, clk, in, r6663_out);
	reg32 r6664 (rst, clk, in, r6664_out);
	reg32 r6665 (rst, clk, in, r6665_out);
	reg32 r6666 (rst, clk, in, r6666_out);
	reg32 r6667 (rst, clk, in, r6667_out);
	reg32 r6668 (rst, clk, in, r6668_out);
	reg32 r6669 (rst, clk, in, r6669_out);
	reg32 r6670 (rst, clk, in, r6670_out);
	reg32 r6671 (rst, clk, in, r6671_out);
	reg32 r6672 (rst, clk, in, r6672_out);
	reg32 r6673 (rst, clk, in, r6673_out);
	reg32 r6674 (rst, clk, in, r6674_out);
	reg32 r6675 (rst, clk, in, r6675_out);
	reg32 r6676 (rst, clk, in, r6676_out);
	reg32 r6677 (rst, clk, in, r6677_out);
	reg32 r6678 (rst, clk, in, r6678_out);
	reg32 r6679 (rst, clk, in, r6679_out);
	reg32 r6680 (rst, clk, in, r6680_out);
	reg32 r6681 (rst, clk, in, r6681_out);
	reg32 r6682 (rst, clk, in, r6682_out);
	reg32 r6683 (rst, clk, in, r6683_out);
	reg32 r6684 (rst, clk, in, r6684_out);
	reg32 r6685 (rst, clk, in, r6685_out);
	reg32 r6686 (rst, clk, in, r6686_out);
	reg32 r6687 (rst, clk, in, r6687_out);
	reg32 r6688 (rst, clk, in, r6688_out);
	reg32 r6689 (rst, clk, in, r6689_out);
	reg32 r6690 (rst, clk, in, r6690_out);
	reg32 r6691 (rst, clk, in, r6691_out);
	reg32 r6692 (rst, clk, in, r6692_out);
	reg32 r6693 (rst, clk, in, r6693_out);
	reg32 r6694 (rst, clk, in, r6694_out);
	reg32 r6695 (rst, clk, in, r6695_out);
	reg32 r6696 (rst, clk, in, r6696_out);
	reg32 r6697 (rst, clk, in, r6697_out);
	reg32 r6698 (rst, clk, in, r6698_out);
	reg32 r6699 (rst, clk, in, r6699_out);
	reg32 r6700 (rst, clk, in, r6700_out);
	reg32 r6701 (rst, clk, in, r6701_out);
	reg32 r6702 (rst, clk, in, r6702_out);
	reg32 r6703 (rst, clk, in, r6703_out);
	reg32 r6704 (rst, clk, in, r6704_out);
	reg32 r6705 (rst, clk, in, r6705_out);
	reg32 r6706 (rst, clk, in, r6706_out);
	reg32 r6707 (rst, clk, in, r6707_out);
	reg32 r6708 (rst, clk, in, r6708_out);
	reg32 r6709 (rst, clk, in, r6709_out);
	reg32 r6710 (rst, clk, in, r6710_out);
	reg32 r6711 (rst, clk, in, r6711_out);
	reg32 r6712 (rst, clk, in, r6712_out);
	reg32 r6713 (rst, clk, in, r6713_out);
	reg32 r6714 (rst, clk, in, r6714_out);
	reg32 r6715 (rst, clk, in, r6715_out);
	reg32 r6716 (rst, clk, in, r6716_out);
	reg32 r6717 (rst, clk, in, r6717_out);
	reg32 r6718 (rst, clk, in, r6718_out);
	reg32 r6719 (rst, clk, in, r6719_out);
	reg32 r6720 (rst, clk, in, r6720_out);
	reg32 r6721 (rst, clk, in, r6721_out);
	reg32 r6722 (rst, clk, in, r6722_out);
	reg32 r6723 (rst, clk, in, r6723_out);
	reg32 r6724 (rst, clk, in, r6724_out);
	reg32 r6725 (rst, clk, in, r6725_out);
	reg32 r6726 (rst, clk, in, r6726_out);
	reg32 r6727 (rst, clk, in, r6727_out);
	reg32 r6728 (rst, clk, in, r6728_out);
	reg32 r6729 (rst, clk, in, r6729_out);
	reg32 r6730 (rst, clk, in, r6730_out);
	reg32 r6731 (rst, clk, in, r6731_out);
	reg32 r6732 (rst, clk, in, r6732_out);
	reg32 r6733 (rst, clk, in, r6733_out);
	reg32 r6734 (rst, clk, in, r6734_out);
	reg32 r6735 (rst, clk, in, r6735_out);
	reg32 r6736 (rst, clk, in, r6736_out);
	reg32 r6737 (rst, clk, in, r6737_out);
	reg32 r6738 (rst, clk, in, r6738_out);
	reg32 r6739 (rst, clk, in, r6739_out);
	reg32 r6740 (rst, clk, in, r6740_out);
	reg32 r6741 (rst, clk, in, r6741_out);
	reg32 r6742 (rst, clk, in, r6742_out);
	reg32 r6743 (rst, clk, in, r6743_out);
	reg32 r6744 (rst, clk, in, r6744_out);
	reg32 r6745 (rst, clk, in, r6745_out);
	reg32 r6746 (rst, clk, in, r6746_out);
	reg32 r6747 (rst, clk, in, r6747_out);
	reg32 r6748 (rst, clk, in, r6748_out);
	reg32 r6749 (rst, clk, in, r6749_out);
	reg32 r6750 (rst, clk, in, r6750_out);
	reg32 r6751 (rst, clk, in, r6751_out);
	reg32 r6752 (rst, clk, in, r6752_out);
	reg32 r6753 (rst, clk, in, r6753_out);
	reg32 r6754 (rst, clk, in, r6754_out);
	reg32 r6755 (rst, clk, in, r6755_out);
	reg32 r6756 (rst, clk, in, r6756_out);
	reg32 r6757 (rst, clk, in, r6757_out);
	reg32 r6758 (rst, clk, in, r6758_out);
	reg32 r6759 (rst, clk, in, r6759_out);
	reg32 r6760 (rst, clk, in, r6760_out);
	reg32 r6761 (rst, clk, in, r6761_out);
	reg32 r6762 (rst, clk, in, r6762_out);
	reg32 r6763 (rst, clk, in, r6763_out);
	reg32 r6764 (rst, clk, in, r6764_out);
	reg32 r6765 (rst, clk, in, r6765_out);
	reg32 r6766 (rst, clk, in, r6766_out);
	reg32 r6767 (rst, clk, in, r6767_out);
	reg32 r6768 (rst, clk, in, r6768_out);
	reg32 r6769 (rst, clk, in, r6769_out);
	reg32 r6770 (rst, clk, in, r6770_out);
	reg32 r6771 (rst, clk, in, r6771_out);
	reg32 r6772 (rst, clk, in, r6772_out);
	reg32 r6773 (rst, clk, in, r6773_out);
	reg32 r6774 (rst, clk, in, r6774_out);
	reg32 r6775 (rst, clk, in, r6775_out);
	reg32 r6776 (rst, clk, in, r6776_out);
	reg32 r6777 (rst, clk, in, r6777_out);
	reg32 r6778 (rst, clk, in, r6778_out);
	reg32 r6779 (rst, clk, in, r6779_out);
	reg32 r6780 (rst, clk, in, r6780_out);
	reg32 r6781 (rst, clk, in, r6781_out);
	reg32 r6782 (rst, clk, in, r6782_out);
	reg32 r6783 (rst, clk, in, r6783_out);
	reg32 r6784 (rst, clk, in, r6784_out);
	reg32 r6785 (rst, clk, in, r6785_out);
	reg32 r6786 (rst, clk, in, r6786_out);
	reg32 r6787 (rst, clk, in, r6787_out);
	reg32 r6788 (rst, clk, in, r6788_out);
	reg32 r6789 (rst, clk, in, r6789_out);
	reg32 r6790 (rst, clk, in, r6790_out);
	reg32 r6791 (rst, clk, in, r6791_out);
	reg32 r6792 (rst, clk, in, r6792_out);
	reg32 r6793 (rst, clk, in, r6793_out);
	reg32 r6794 (rst, clk, in, r6794_out);
	reg32 r6795 (rst, clk, in, r6795_out);
	reg32 r6796 (rst, clk, in, r6796_out);
	reg32 r6797 (rst, clk, in, r6797_out);
	reg32 r6798 (rst, clk, in, r6798_out);
	reg32 r6799 (rst, clk, in, r6799_out);
	reg32 r6800 (rst, clk, in, r6800_out);
	reg32 r6801 (rst, clk, in, r6801_out);
	reg32 r6802 (rst, clk, in, r6802_out);
	reg32 r6803 (rst, clk, in, r6803_out);
	reg32 r6804 (rst, clk, in, r6804_out);
	reg32 r6805 (rst, clk, in, r6805_out);
	reg32 r6806 (rst, clk, in, r6806_out);
	reg32 r6807 (rst, clk, in, r6807_out);
	reg32 r6808 (rst, clk, in, r6808_out);
	reg32 r6809 (rst, clk, in, r6809_out);
	reg32 r6810 (rst, clk, in, r6810_out);
	reg32 r6811 (rst, clk, in, r6811_out);
	reg32 r6812 (rst, clk, in, r6812_out);
	reg32 r6813 (rst, clk, in, r6813_out);
	reg32 r6814 (rst, clk, in, r6814_out);
	reg32 r6815 (rst, clk, in, r6815_out);
	reg32 r6816 (rst, clk, in, r6816_out);
	reg32 r6817 (rst, clk, in, r6817_out);
	reg32 r6818 (rst, clk, in, r6818_out);
	reg32 r6819 (rst, clk, in, r6819_out);
	reg32 r6820 (rst, clk, in, r6820_out);
	reg32 r6821 (rst, clk, in, r6821_out);
	reg32 r6822 (rst, clk, in, r6822_out);
	reg32 r6823 (rst, clk, in, r6823_out);
	reg32 r6824 (rst, clk, in, r6824_out);
	reg32 r6825 (rst, clk, in, r6825_out);
	reg32 r6826 (rst, clk, in, r6826_out);
	reg32 r6827 (rst, clk, in, r6827_out);
	reg32 r6828 (rst, clk, in, r6828_out);
	reg32 r6829 (rst, clk, in, r6829_out);
	reg32 r6830 (rst, clk, in, r6830_out);
	reg32 r6831 (rst, clk, in, r6831_out);
	reg32 r6832 (rst, clk, in, r6832_out);
	reg32 r6833 (rst, clk, in, r6833_out);
	reg32 r6834 (rst, clk, in, r6834_out);
	reg32 r6835 (rst, clk, in, r6835_out);
	reg32 r6836 (rst, clk, in, r6836_out);
	reg32 r6837 (rst, clk, in, r6837_out);
	reg32 r6838 (rst, clk, in, r6838_out);
	reg32 r6839 (rst, clk, in, r6839_out);
	reg32 r6840 (rst, clk, in, r6840_out);
	reg32 r6841 (rst, clk, in, r6841_out);
	reg32 r6842 (rst, clk, in, r6842_out);
	reg32 r6843 (rst, clk, in, r6843_out);
	reg32 r6844 (rst, clk, in, r6844_out);
	reg32 r6845 (rst, clk, in, r6845_out);
	reg32 r6846 (rst, clk, in, r6846_out);
	reg32 r6847 (rst, clk, in, r6847_out);
	reg32 r6848 (rst, clk, in, r6848_out);
	reg32 r6849 (rst, clk, in, r6849_out);
	reg32 r6850 (rst, clk, in, r6850_out);
	reg32 r6851 (rst, clk, in, r6851_out);
	reg32 r6852 (rst, clk, in, r6852_out);
	reg32 r6853 (rst, clk, in, r6853_out);
	reg32 r6854 (rst, clk, in, r6854_out);
	reg32 r6855 (rst, clk, in, r6855_out);
	reg32 r6856 (rst, clk, in, r6856_out);
	reg32 r6857 (rst, clk, in, r6857_out);
	reg32 r6858 (rst, clk, in, r6858_out);
	reg32 r6859 (rst, clk, in, r6859_out);
	reg32 r6860 (rst, clk, in, r6860_out);
	reg32 r6861 (rst, clk, in, r6861_out);
	reg32 r6862 (rst, clk, in, r6862_out);
	reg32 r6863 (rst, clk, in, r6863_out);
	reg32 r6864 (rst, clk, in, r6864_out);
	reg32 r6865 (rst, clk, in, r6865_out);
	reg32 r6866 (rst, clk, in, r6866_out);
	reg32 r6867 (rst, clk, in, r6867_out);
	reg32 r6868 (rst, clk, in, r6868_out);
	reg32 r6869 (rst, clk, in, r6869_out);
	reg32 r6870 (rst, clk, in, r6870_out);
	reg32 r6871 (rst, clk, in, r6871_out);
	reg32 r6872 (rst, clk, in, r6872_out);
	reg32 r6873 (rst, clk, in, r6873_out);
	reg32 r6874 (rst, clk, in, r6874_out);
	reg32 r6875 (rst, clk, in, r6875_out);
	reg32 r6876 (rst, clk, in, r6876_out);
	reg32 r6877 (rst, clk, in, r6877_out);
	reg32 r6878 (rst, clk, in, r6878_out);
	reg32 r6879 (rst, clk, in, r6879_out);
	reg32 r6880 (rst, clk, in, r6880_out);
	reg32 r6881 (rst, clk, in, r6881_out);
	reg32 r6882 (rst, clk, in, r6882_out);
	reg32 r6883 (rst, clk, in, r6883_out);
	reg32 r6884 (rst, clk, in, r6884_out);
	reg32 r6885 (rst, clk, in, r6885_out);
	reg32 r6886 (rst, clk, in, r6886_out);
	reg32 r6887 (rst, clk, in, r6887_out);
	reg32 r6888 (rst, clk, in, r6888_out);
	reg32 r6889 (rst, clk, in, r6889_out);
	reg32 r6890 (rst, clk, in, r6890_out);
	reg32 r6891 (rst, clk, in, r6891_out);
	reg32 r6892 (rst, clk, in, r6892_out);
	reg32 r6893 (rst, clk, in, r6893_out);
	reg32 r6894 (rst, clk, in, r6894_out);
	reg32 r6895 (rst, clk, in, r6895_out);
	reg32 r6896 (rst, clk, in, r6896_out);
	reg32 r6897 (rst, clk, in, r6897_out);
	reg32 r6898 (rst, clk, in, r6898_out);
	reg32 r6899 (rst, clk, in, r6899_out);
	reg32 r6900 (rst, clk, in, r6900_out);
	reg32 r6901 (rst, clk, in, r6901_out);
	reg32 r6902 (rst, clk, in, r6902_out);
	reg32 r6903 (rst, clk, in, r6903_out);
	reg32 r6904 (rst, clk, in, r6904_out);
	reg32 r6905 (rst, clk, in, r6905_out);
	reg32 r6906 (rst, clk, in, r6906_out);
	reg32 r6907 (rst, clk, in, r6907_out);
	reg32 r6908 (rst, clk, in, r6908_out);
	reg32 r6909 (rst, clk, in, r6909_out);
	reg32 r6910 (rst, clk, in, r6910_out);
	reg32 r6911 (rst, clk, in, r6911_out);
	reg32 r6912 (rst, clk, in, r6912_out);
	reg32 r6913 (rst, clk, in, r6913_out);
	reg32 r6914 (rst, clk, in, r6914_out);
	reg32 r6915 (rst, clk, in, r6915_out);
	reg32 r6916 (rst, clk, in, r6916_out);
	reg32 r6917 (rst, clk, in, r6917_out);
	reg32 r6918 (rst, clk, in, r6918_out);
	reg32 r6919 (rst, clk, in, r6919_out);
	reg32 r6920 (rst, clk, in, r6920_out);
	reg32 r6921 (rst, clk, in, r6921_out);
	reg32 r6922 (rst, clk, in, r6922_out);
	reg32 r6923 (rst, clk, in, r6923_out);
	reg32 r6924 (rst, clk, in, r6924_out);
	reg32 r6925 (rst, clk, in, r6925_out);
	reg32 r6926 (rst, clk, in, r6926_out);
	reg32 r6927 (rst, clk, in, r6927_out);
	reg32 r6928 (rst, clk, in, r6928_out);
	reg32 r6929 (rst, clk, in, r6929_out);
	reg32 r6930 (rst, clk, in, r6930_out);
	reg32 r6931 (rst, clk, in, r6931_out);
	reg32 r6932 (rst, clk, in, r6932_out);
	reg32 r6933 (rst, clk, in, r6933_out);
	reg32 r6934 (rst, clk, in, r6934_out);
	reg32 r6935 (rst, clk, in, r6935_out);
	reg32 r6936 (rst, clk, in, r6936_out);
	reg32 r6937 (rst, clk, in, r6937_out);
	reg32 r6938 (rst, clk, in, r6938_out);
	reg32 r6939 (rst, clk, in, r6939_out);
	reg32 r6940 (rst, clk, in, r6940_out);
	reg32 r6941 (rst, clk, in, r6941_out);
	reg32 r6942 (rst, clk, in, r6942_out);
	reg32 r6943 (rst, clk, in, r6943_out);
	reg32 r6944 (rst, clk, in, r6944_out);
	reg32 r6945 (rst, clk, in, r6945_out);
	reg32 r6946 (rst, clk, in, r6946_out);
	reg32 r6947 (rst, clk, in, r6947_out);
	reg32 r6948 (rst, clk, in, r6948_out);
	reg32 r6949 (rst, clk, in, r6949_out);
	reg32 r6950 (rst, clk, in, r6950_out);
	reg32 r6951 (rst, clk, in, r6951_out);
	reg32 r6952 (rst, clk, in, r6952_out);
	reg32 r6953 (rst, clk, in, r6953_out);
	reg32 r6954 (rst, clk, in, r6954_out);
	reg32 r6955 (rst, clk, in, r6955_out);
	reg32 r6956 (rst, clk, in, r6956_out);
	reg32 r6957 (rst, clk, in, r6957_out);
	reg32 r6958 (rst, clk, in, r6958_out);
	reg32 r6959 (rst, clk, in, r6959_out);
	reg32 r6960 (rst, clk, in, r6960_out);
	reg32 r6961 (rst, clk, in, r6961_out);
	reg32 r6962 (rst, clk, in, r6962_out);
	reg32 r6963 (rst, clk, in, r6963_out);
	reg32 r6964 (rst, clk, in, r6964_out);
	reg32 r6965 (rst, clk, in, r6965_out);
	reg32 r6966 (rst, clk, in, r6966_out);
	reg32 r6967 (rst, clk, in, r6967_out);
	reg32 r6968 (rst, clk, in, r6968_out);
	reg32 r6969 (rst, clk, in, r6969_out);
	reg32 r6970 (rst, clk, in, r6970_out);
	reg32 r6971 (rst, clk, in, r6971_out);
	reg32 r6972 (rst, clk, in, r6972_out);
	reg32 r6973 (rst, clk, in, r6973_out);
	reg32 r6974 (rst, clk, in, r6974_out);
	reg32 r6975 (rst, clk, in, r6975_out);
	reg32 r6976 (rst, clk, in, r6976_out);
	reg32 r6977 (rst, clk, in, r6977_out);
	reg32 r6978 (rst, clk, in, r6978_out);
	reg32 r6979 (rst, clk, in, r6979_out);
	reg32 r6980 (rst, clk, in, r6980_out);
	reg32 r6981 (rst, clk, in, r6981_out);
	reg32 r6982 (rst, clk, in, r6982_out);
	reg32 r6983 (rst, clk, in, r6983_out);
	reg32 r6984 (rst, clk, in, r6984_out);
	reg32 r6985 (rst, clk, in, r6985_out);
	reg32 r6986 (rst, clk, in, r6986_out);
	reg32 r6987 (rst, clk, in, r6987_out);
	reg32 r6988 (rst, clk, in, r6988_out);
	reg32 r6989 (rst, clk, in, r6989_out);
	reg32 r6990 (rst, clk, in, r6990_out);
	reg32 r6991 (rst, clk, in, r6991_out);
	reg32 r6992 (rst, clk, in, r6992_out);
	reg32 r6993 (rst, clk, in, r6993_out);
	reg32 r6994 (rst, clk, in, r6994_out);
	reg32 r6995 (rst, clk, in, r6995_out);
	reg32 r6996 (rst, clk, in, r6996_out);
	reg32 r6997 (rst, clk, in, r6997_out);
	reg32 r6998 (rst, clk, in, r6998_out);
	reg32 r6999 (rst, clk, in, r6999_out);
	reg32 r7000 (rst, clk, in, r7000_out);
	reg32 r7001 (rst, clk, in, r7001_out);
	reg32 r7002 (rst, clk, in, r7002_out);
	reg32 r7003 (rst, clk, in, r7003_out);
	reg32 r7004 (rst, clk, in, r7004_out);
	reg32 r7005 (rst, clk, in, r7005_out);
	reg32 r7006 (rst, clk, in, r7006_out);
	reg32 r7007 (rst, clk, in, r7007_out);
	reg32 r7008 (rst, clk, in, r7008_out);
	reg32 r7009 (rst, clk, in, r7009_out);
	reg32 r7010 (rst, clk, in, r7010_out);
	reg32 r7011 (rst, clk, in, r7011_out);
	reg32 r7012 (rst, clk, in, r7012_out);
	reg32 r7013 (rst, clk, in, r7013_out);
	reg32 r7014 (rst, clk, in, r7014_out);
	reg32 r7015 (rst, clk, in, r7015_out);
	reg32 r7016 (rst, clk, in, r7016_out);
	reg32 r7017 (rst, clk, in, r7017_out);
	reg32 r7018 (rst, clk, in, r7018_out);
	reg32 r7019 (rst, clk, in, r7019_out);
	reg32 r7020 (rst, clk, in, r7020_out);
	reg32 r7021 (rst, clk, in, r7021_out);
	reg32 r7022 (rst, clk, in, r7022_out);
	reg32 r7023 (rst, clk, in, r7023_out);
	reg32 r7024 (rst, clk, in, r7024_out);
	reg32 r7025 (rst, clk, in, r7025_out);
	reg32 r7026 (rst, clk, in, r7026_out);
	reg32 r7027 (rst, clk, in, r7027_out);
	reg32 r7028 (rst, clk, in, r7028_out);
	reg32 r7029 (rst, clk, in, r7029_out);
	reg32 r7030 (rst, clk, in, r7030_out);
	reg32 r7031 (rst, clk, in, r7031_out);
	reg32 r7032 (rst, clk, in, r7032_out);
	reg32 r7033 (rst, clk, in, r7033_out);
	reg32 r7034 (rst, clk, in, r7034_out);
	reg32 r7035 (rst, clk, in, r7035_out);
	reg32 r7036 (rst, clk, in, r7036_out);
	reg32 r7037 (rst, clk, in, r7037_out);
	reg32 r7038 (rst, clk, in, r7038_out);
	reg32 r7039 (rst, clk, in, r7039_out);
	reg32 r7040 (rst, clk, in, r7040_out);
	reg32 r7041 (rst, clk, in, r7041_out);
	reg32 r7042 (rst, clk, in, r7042_out);
	reg32 r7043 (rst, clk, in, r7043_out);
	reg32 r7044 (rst, clk, in, r7044_out);
	reg32 r7045 (rst, clk, in, r7045_out);
	reg32 r7046 (rst, clk, in, r7046_out);
	reg32 r7047 (rst, clk, in, r7047_out);
	reg32 r7048 (rst, clk, in, r7048_out);
	reg32 r7049 (rst, clk, in, r7049_out);
	reg32 r7050 (rst, clk, in, r7050_out);
	reg32 r7051 (rst, clk, in, r7051_out);
	reg32 r7052 (rst, clk, in, r7052_out);
	reg32 r7053 (rst, clk, in, r7053_out);
	reg32 r7054 (rst, clk, in, r7054_out);
	reg32 r7055 (rst, clk, in, r7055_out);
	reg32 r7056 (rst, clk, in, r7056_out);
	reg32 r7057 (rst, clk, in, r7057_out);
	reg32 r7058 (rst, clk, in, r7058_out);
	reg32 r7059 (rst, clk, in, r7059_out);
	reg32 r7060 (rst, clk, in, r7060_out);
	reg32 r7061 (rst, clk, in, r7061_out);
	reg32 r7062 (rst, clk, in, r7062_out);
	reg32 r7063 (rst, clk, in, r7063_out);
	reg32 r7064 (rst, clk, in, r7064_out);
	reg32 r7065 (rst, clk, in, r7065_out);
	reg32 r7066 (rst, clk, in, r7066_out);
	reg32 r7067 (rst, clk, in, r7067_out);
	reg32 r7068 (rst, clk, in, r7068_out);
	reg32 r7069 (rst, clk, in, r7069_out);
	reg32 r7070 (rst, clk, in, r7070_out);
	reg32 r7071 (rst, clk, in, r7071_out);
	reg32 r7072 (rst, clk, in, r7072_out);
	reg32 r7073 (rst, clk, in, r7073_out);
	reg32 r7074 (rst, clk, in, r7074_out);
	reg32 r7075 (rst, clk, in, r7075_out);
	reg32 r7076 (rst, clk, in, r7076_out);
	reg32 r7077 (rst, clk, in, r7077_out);
	reg32 r7078 (rst, clk, in, r7078_out);
	reg32 r7079 (rst, clk, in, r7079_out);
	reg32 r7080 (rst, clk, in, r7080_out);
	reg32 r7081 (rst, clk, in, r7081_out);
	reg32 r7082 (rst, clk, in, r7082_out);
	reg32 r7083 (rst, clk, in, r7083_out);
	reg32 r7084 (rst, clk, in, r7084_out);
	reg32 r7085 (rst, clk, in, r7085_out);
	reg32 r7086 (rst, clk, in, r7086_out);
	reg32 r7087 (rst, clk, in, r7087_out);
	reg32 r7088 (rst, clk, in, r7088_out);
	reg32 r7089 (rst, clk, in, r7089_out);
	reg32 r7090 (rst, clk, in, r7090_out);
	reg32 r7091 (rst, clk, in, r7091_out);
	reg32 r7092 (rst, clk, in, r7092_out);
	reg32 r7093 (rst, clk, in, r7093_out);
	reg32 r7094 (rst, clk, in, r7094_out);
	reg32 r7095 (rst, clk, in, r7095_out);
	reg32 r7096 (rst, clk, in, r7096_out);
	reg32 r7097 (rst, clk, in, r7097_out);
	reg32 r7098 (rst, clk, in, r7098_out);
	reg32 r7099 (rst, clk, in, r7099_out);
	reg32 r7100 (rst, clk, in, r7100_out);
	reg32 r7101 (rst, clk, in, r7101_out);
	reg32 r7102 (rst, clk, in, r7102_out);
	reg32 r7103 (rst, clk, in, r7103_out);
	reg32 r7104 (rst, clk, in, r7104_out);
	reg32 r7105 (rst, clk, in, r7105_out);
	reg32 r7106 (rst, clk, in, r7106_out);
	reg32 r7107 (rst, clk, in, r7107_out);
	reg32 r7108 (rst, clk, in, r7108_out);
	reg32 r7109 (rst, clk, in, r7109_out);
	reg32 r7110 (rst, clk, in, r7110_out);
	reg32 r7111 (rst, clk, in, r7111_out);
	reg32 r7112 (rst, clk, in, r7112_out);
	reg32 r7113 (rst, clk, in, r7113_out);
	reg32 r7114 (rst, clk, in, r7114_out);
	reg32 r7115 (rst, clk, in, r7115_out);
	reg32 r7116 (rst, clk, in, r7116_out);
	reg32 r7117 (rst, clk, in, r7117_out);
	reg32 r7118 (rst, clk, in, r7118_out);
	reg32 r7119 (rst, clk, in, r7119_out);
	reg32 r7120 (rst, clk, in, r7120_out);
	reg32 r7121 (rst, clk, in, r7121_out);
	reg32 r7122 (rst, clk, in, r7122_out);
	reg32 r7123 (rst, clk, in, r7123_out);
	reg32 r7124 (rst, clk, in, r7124_out);
	reg32 r7125 (rst, clk, in, r7125_out);
	reg32 r7126 (rst, clk, in, r7126_out);
	reg32 r7127 (rst, clk, in, r7127_out);
	reg32 r7128 (rst, clk, in, r7128_out);
	reg32 r7129 (rst, clk, in, r7129_out);
	reg32 r7130 (rst, clk, in, r7130_out);
	reg32 r7131 (rst, clk, in, r7131_out);
	reg32 r7132 (rst, clk, in, r7132_out);
	reg32 r7133 (rst, clk, in, r7133_out);
	reg32 r7134 (rst, clk, in, r7134_out);
	reg32 r7135 (rst, clk, in, r7135_out);
	reg32 r7136 (rst, clk, in, r7136_out);
	reg32 r7137 (rst, clk, in, r7137_out);
	reg32 r7138 (rst, clk, in, r7138_out);
	reg32 r7139 (rst, clk, in, r7139_out);
	reg32 r7140 (rst, clk, in, r7140_out);
	reg32 r7141 (rst, clk, in, r7141_out);
	reg32 r7142 (rst, clk, in, r7142_out);
	reg32 r7143 (rst, clk, in, r7143_out);
	reg32 r7144 (rst, clk, in, r7144_out);
	reg32 r7145 (rst, clk, in, r7145_out);
	reg32 r7146 (rst, clk, in, r7146_out);
	reg32 r7147 (rst, clk, in, r7147_out);
	reg32 r7148 (rst, clk, in, r7148_out);
	reg32 r7149 (rst, clk, in, r7149_out);
	reg32 r7150 (rst, clk, in, r7150_out);
	reg32 r7151 (rst, clk, in, r7151_out);
	reg32 r7152 (rst, clk, in, r7152_out);
	reg32 r7153 (rst, clk, in, r7153_out);
	reg32 r7154 (rst, clk, in, r7154_out);
	reg32 r7155 (rst, clk, in, r7155_out);
	reg32 r7156 (rst, clk, in, r7156_out);
	reg32 r7157 (rst, clk, in, r7157_out);
	reg32 r7158 (rst, clk, in, r7158_out);
	reg32 r7159 (rst, clk, in, r7159_out);
	reg32 r7160 (rst, clk, in, r7160_out);
	reg32 r7161 (rst, clk, in, r7161_out);
	reg32 r7162 (rst, clk, in, r7162_out);
	reg32 r7163 (rst, clk, in, r7163_out);
	reg32 r7164 (rst, clk, in, r7164_out);
	reg32 r7165 (rst, clk, in, r7165_out);
	reg32 r7166 (rst, clk, in, r7166_out);
	reg32 r7167 (rst, clk, in, r7167_out);
	reg32 r7168 (rst, clk, in, r7168_out);
	reg32 r7169 (rst, clk, in, r7169_out);
	reg32 r7170 (rst, clk, in, r7170_out);
	reg32 r7171 (rst, clk, in, r7171_out);
	reg32 r7172 (rst, clk, in, r7172_out);
	reg32 r7173 (rst, clk, in, r7173_out);
	reg32 r7174 (rst, clk, in, r7174_out);
	reg32 r7175 (rst, clk, in, r7175_out);
	reg32 r7176 (rst, clk, in, r7176_out);
	reg32 r7177 (rst, clk, in, r7177_out);
	reg32 r7178 (rst, clk, in, r7178_out);
	reg32 r7179 (rst, clk, in, r7179_out);
	reg32 r7180 (rst, clk, in, r7180_out);
	reg32 r7181 (rst, clk, in, r7181_out);
	reg32 r7182 (rst, clk, in, r7182_out);
	reg32 r7183 (rst, clk, in, r7183_out);
	reg32 r7184 (rst, clk, in, r7184_out);
	reg32 r7185 (rst, clk, in, r7185_out);
	reg32 r7186 (rst, clk, in, r7186_out);
	reg32 r7187 (rst, clk, in, r7187_out);
	reg32 r7188 (rst, clk, in, r7188_out);
	reg32 r7189 (rst, clk, in, r7189_out);
	reg32 r7190 (rst, clk, in, r7190_out);
	reg32 r7191 (rst, clk, in, r7191_out);
	reg32 r7192 (rst, clk, in, r7192_out);
	reg32 r7193 (rst, clk, in, r7193_out);
	reg32 r7194 (rst, clk, in, r7194_out);
	reg32 r7195 (rst, clk, in, r7195_out);
	reg32 r7196 (rst, clk, in, r7196_out);
	reg32 r7197 (rst, clk, in, r7197_out);
	reg32 r7198 (rst, clk, in, r7198_out);
	reg32 r7199 (rst, clk, in, r7199_out);
	reg32 r7200 (rst, clk, in, r7200_out);
	reg32 r7201 (rst, clk, in, r7201_out);
	reg32 r7202 (rst, clk, in, r7202_out);
	reg32 r7203 (rst, clk, in, r7203_out);
	reg32 r7204 (rst, clk, in, r7204_out);
	reg32 r7205 (rst, clk, in, r7205_out);
	reg32 r7206 (rst, clk, in, r7206_out);
	reg32 r7207 (rst, clk, in, r7207_out);
	reg32 r7208 (rst, clk, in, r7208_out);
	reg32 r7209 (rst, clk, in, r7209_out);
	reg32 r7210 (rst, clk, in, r7210_out);
	reg32 r7211 (rst, clk, in, r7211_out);
	reg32 r7212 (rst, clk, in, r7212_out);
	reg32 r7213 (rst, clk, in, r7213_out);
	reg32 r7214 (rst, clk, in, r7214_out);
	reg32 r7215 (rst, clk, in, r7215_out);
	reg32 r7216 (rst, clk, in, r7216_out);
	reg32 r7217 (rst, clk, in, r7217_out);
	reg32 r7218 (rst, clk, in, r7218_out);
	reg32 r7219 (rst, clk, in, r7219_out);
	reg32 r7220 (rst, clk, in, r7220_out);
	reg32 r7221 (rst, clk, in, r7221_out);
	reg32 r7222 (rst, clk, in, r7222_out);
	reg32 r7223 (rst, clk, in, r7223_out);
	reg32 r7224 (rst, clk, in, r7224_out);
	reg32 r7225 (rst, clk, in, r7225_out);
	reg32 r7226 (rst, clk, in, r7226_out);
	reg32 r7227 (rst, clk, in, r7227_out);
	reg32 r7228 (rst, clk, in, r7228_out);
	reg32 r7229 (rst, clk, in, r7229_out);
	reg32 r7230 (rst, clk, in, r7230_out);
	reg32 r7231 (rst, clk, in, r7231_out);
	reg32 r7232 (rst, clk, in, r7232_out);
	reg32 r7233 (rst, clk, in, r7233_out);
	reg32 r7234 (rst, clk, in, r7234_out);
	reg32 r7235 (rst, clk, in, r7235_out);
	reg32 r7236 (rst, clk, in, r7236_out);
	reg32 r7237 (rst, clk, in, r7237_out);
	reg32 r7238 (rst, clk, in, r7238_out);
	reg32 r7239 (rst, clk, in, r7239_out);
	reg32 r7240 (rst, clk, in, r7240_out);
	reg32 r7241 (rst, clk, in, r7241_out);
	reg32 r7242 (rst, clk, in, r7242_out);
	reg32 r7243 (rst, clk, in, r7243_out);
	reg32 r7244 (rst, clk, in, r7244_out);
	reg32 r7245 (rst, clk, in, r7245_out);
	reg32 r7246 (rst, clk, in, r7246_out);
	reg32 r7247 (rst, clk, in, r7247_out);
	reg32 r7248 (rst, clk, in, r7248_out);
	reg32 r7249 (rst, clk, in, r7249_out);
	reg32 r7250 (rst, clk, in, r7250_out);
	reg32 r7251 (rst, clk, in, r7251_out);
	reg32 r7252 (rst, clk, in, r7252_out);
	reg32 r7253 (rst, clk, in, r7253_out);
	reg32 r7254 (rst, clk, in, r7254_out);
	reg32 r7255 (rst, clk, in, r7255_out);
	reg32 r7256 (rst, clk, in, r7256_out);
	reg32 r7257 (rst, clk, in, r7257_out);
	reg32 r7258 (rst, clk, in, r7258_out);
	reg32 r7259 (rst, clk, in, r7259_out);
	reg32 r7260 (rst, clk, in, r7260_out);
	reg32 r7261 (rst, clk, in, r7261_out);
	reg32 r7262 (rst, clk, in, r7262_out);
	reg32 r7263 (rst, clk, in, r7263_out);
	reg32 r7264 (rst, clk, in, r7264_out);
	reg32 r7265 (rst, clk, in, r7265_out);
	reg32 r7266 (rst, clk, in, r7266_out);
	reg32 r7267 (rst, clk, in, r7267_out);
	reg32 r7268 (rst, clk, in, r7268_out);
	reg32 r7269 (rst, clk, in, r7269_out);
	reg32 r7270 (rst, clk, in, r7270_out);
	reg32 r7271 (rst, clk, in, r7271_out);
	reg32 r7272 (rst, clk, in, r7272_out);
	reg32 r7273 (rst, clk, in, r7273_out);
	reg32 r7274 (rst, clk, in, r7274_out);
	reg32 r7275 (rst, clk, in, r7275_out);
	reg32 r7276 (rst, clk, in, r7276_out);
	reg32 r7277 (rst, clk, in, r7277_out);
	reg32 r7278 (rst, clk, in, r7278_out);
	reg32 r7279 (rst, clk, in, r7279_out);
	reg32 r7280 (rst, clk, in, r7280_out);
	reg32 r7281 (rst, clk, in, r7281_out);
	reg32 r7282 (rst, clk, in, r7282_out);
	reg32 r7283 (rst, clk, in, r7283_out);
	reg32 r7284 (rst, clk, in, r7284_out);
	reg32 r7285 (rst, clk, in, r7285_out);
	reg32 r7286 (rst, clk, in, r7286_out);
	reg32 r7287 (rst, clk, in, r7287_out);
	reg32 r7288 (rst, clk, in, r7288_out);
	reg32 r7289 (rst, clk, in, r7289_out);
	reg32 r7290 (rst, clk, in, r7290_out);
	reg32 r7291 (rst, clk, in, r7291_out);
	reg32 r7292 (rst, clk, in, r7292_out);
	reg32 r7293 (rst, clk, in, r7293_out);
	reg32 r7294 (rst, clk, in, r7294_out);
	reg32 r7295 (rst, clk, in, r7295_out);
	reg32 r7296 (rst, clk, in, r7296_out);
	reg32 r7297 (rst, clk, in, r7297_out);
	reg32 r7298 (rst, clk, in, r7298_out);
	reg32 r7299 (rst, clk, in, r7299_out);
	reg32 r7300 (rst, clk, in, r7300_out);
	reg32 r7301 (rst, clk, in, r7301_out);
	reg32 r7302 (rst, clk, in, r7302_out);
	reg32 r7303 (rst, clk, in, r7303_out);
	reg32 r7304 (rst, clk, in, r7304_out);
	reg32 r7305 (rst, clk, in, r7305_out);
	reg32 r7306 (rst, clk, in, r7306_out);
	reg32 r7307 (rst, clk, in, r7307_out);
	reg32 r7308 (rst, clk, in, r7308_out);
	reg32 r7309 (rst, clk, in, r7309_out);
	reg32 r7310 (rst, clk, in, r7310_out);
	reg32 r7311 (rst, clk, in, r7311_out);
	reg32 r7312 (rst, clk, in, r7312_out);
	reg32 r7313 (rst, clk, in, r7313_out);
	reg32 r7314 (rst, clk, in, r7314_out);
	reg32 r7315 (rst, clk, in, r7315_out);
	reg32 r7316 (rst, clk, in, r7316_out);
	reg32 r7317 (rst, clk, in, r7317_out);
	reg32 r7318 (rst, clk, in, r7318_out);
	reg32 r7319 (rst, clk, in, r7319_out);
	reg32 r7320 (rst, clk, in, r7320_out);
	reg32 r7321 (rst, clk, in, r7321_out);
	reg32 r7322 (rst, clk, in, r7322_out);
	reg32 r7323 (rst, clk, in, r7323_out);
	reg32 r7324 (rst, clk, in, r7324_out);
	reg32 r7325 (rst, clk, in, r7325_out);
	reg32 r7326 (rst, clk, in, r7326_out);
	reg32 r7327 (rst, clk, in, r7327_out);
	reg32 r7328 (rst, clk, in, r7328_out);
	reg32 r7329 (rst, clk, in, r7329_out);
	reg32 r7330 (rst, clk, in, r7330_out);
	reg32 r7331 (rst, clk, in, r7331_out);
	reg32 r7332 (rst, clk, in, r7332_out);
	reg32 r7333 (rst, clk, in, r7333_out);
	reg32 r7334 (rst, clk, in, r7334_out);
	reg32 r7335 (rst, clk, in, r7335_out);
	reg32 r7336 (rst, clk, in, r7336_out);
	reg32 r7337 (rst, clk, in, r7337_out);
	reg32 r7338 (rst, clk, in, r7338_out);
	reg32 r7339 (rst, clk, in, r7339_out);
	reg32 r7340 (rst, clk, in, r7340_out);
	reg32 r7341 (rst, clk, in, r7341_out);
	reg32 r7342 (rst, clk, in, r7342_out);
	reg32 r7343 (rst, clk, in, r7343_out);
	reg32 r7344 (rst, clk, in, r7344_out);
	reg32 r7345 (rst, clk, in, r7345_out);
	reg32 r7346 (rst, clk, in, r7346_out);
	reg32 r7347 (rst, clk, in, r7347_out);
	reg32 r7348 (rst, clk, in, r7348_out);
	reg32 r7349 (rst, clk, in, r7349_out);
	reg32 r7350 (rst, clk, in, r7350_out);
	reg32 r7351 (rst, clk, in, r7351_out);
	reg32 r7352 (rst, clk, in, r7352_out);
	reg32 r7353 (rst, clk, in, r7353_out);
	reg32 r7354 (rst, clk, in, r7354_out);
	reg32 r7355 (rst, clk, in, r7355_out);
	reg32 r7356 (rst, clk, in, r7356_out);
	reg32 r7357 (rst, clk, in, r7357_out);
	reg32 r7358 (rst, clk, in, r7358_out);
	reg32 r7359 (rst, clk, in, r7359_out);
	reg32 r7360 (rst, clk, in, r7360_out);
	reg32 r7361 (rst, clk, in, r7361_out);
	reg32 r7362 (rst, clk, in, r7362_out);
	reg32 r7363 (rst, clk, in, r7363_out);
	reg32 r7364 (rst, clk, in, r7364_out);
	reg32 r7365 (rst, clk, in, r7365_out);
	reg32 r7366 (rst, clk, in, r7366_out);
	reg32 r7367 (rst, clk, in, r7367_out);
	reg32 r7368 (rst, clk, in, r7368_out);
	reg32 r7369 (rst, clk, in, r7369_out);
	reg32 r7370 (rst, clk, in, r7370_out);
	reg32 r7371 (rst, clk, in, r7371_out);
	reg32 r7372 (rst, clk, in, r7372_out);
	reg32 r7373 (rst, clk, in, r7373_out);
	reg32 r7374 (rst, clk, in, r7374_out);
	reg32 r7375 (rst, clk, in, r7375_out);
	reg32 r7376 (rst, clk, in, r7376_out);
	reg32 r7377 (rst, clk, in, r7377_out);
	reg32 r7378 (rst, clk, in, r7378_out);
	reg32 r7379 (rst, clk, in, r7379_out);
	reg32 r7380 (rst, clk, in, r7380_out);
	reg32 r7381 (rst, clk, in, r7381_out);
	reg32 r7382 (rst, clk, in, r7382_out);
	reg32 r7383 (rst, clk, in, r7383_out);
	reg32 r7384 (rst, clk, in, r7384_out);
	reg32 r7385 (rst, clk, in, r7385_out);
	reg32 r7386 (rst, clk, in, r7386_out);
	reg32 r7387 (rst, clk, in, r7387_out);
	reg32 r7388 (rst, clk, in, r7388_out);
	reg32 r7389 (rst, clk, in, r7389_out);
	reg32 r7390 (rst, clk, in, r7390_out);
	reg32 r7391 (rst, clk, in, r7391_out);
	reg32 r7392 (rst, clk, in, r7392_out);
	reg32 r7393 (rst, clk, in, r7393_out);
	reg32 r7394 (rst, clk, in, r7394_out);
	reg32 r7395 (rst, clk, in, r7395_out);
	reg32 r7396 (rst, clk, in, r7396_out);
	reg32 r7397 (rst, clk, in, r7397_out);
	reg32 r7398 (rst, clk, in, r7398_out);
	reg32 r7399 (rst, clk, in, r7399_out);
	reg32 r7400 (rst, clk, in, r7400_out);
	reg32 r7401 (rst, clk, in, r7401_out);
	reg32 r7402 (rst, clk, in, r7402_out);
	reg32 r7403 (rst, clk, in, r7403_out);
	reg32 r7404 (rst, clk, in, r7404_out);
	reg32 r7405 (rst, clk, in, r7405_out);
	reg32 r7406 (rst, clk, in, r7406_out);
	reg32 r7407 (rst, clk, in, r7407_out);
	reg32 r7408 (rst, clk, in, r7408_out);
	reg32 r7409 (rst, clk, in, r7409_out);
	reg32 r7410 (rst, clk, in, r7410_out);
	reg32 r7411 (rst, clk, in, r7411_out);
	reg32 r7412 (rst, clk, in, r7412_out);
	reg32 r7413 (rst, clk, in, r7413_out);
	reg32 r7414 (rst, clk, in, r7414_out);
	reg32 r7415 (rst, clk, in, r7415_out);
	reg32 r7416 (rst, clk, in, r7416_out);
	reg32 r7417 (rst, clk, in, r7417_out);
	reg32 r7418 (rst, clk, in, r7418_out);
	reg32 r7419 (rst, clk, in, r7419_out);
	reg32 r7420 (rst, clk, in, r7420_out);
	reg32 r7421 (rst, clk, in, r7421_out);
	reg32 r7422 (rst, clk, in, r7422_out);
	reg32 r7423 (rst, clk, in, r7423_out);
	reg32 r7424 (rst, clk, in, r7424_out);
	reg32 r7425 (rst, clk, in, r7425_out);
	reg32 r7426 (rst, clk, in, r7426_out);
	reg32 r7427 (rst, clk, in, r7427_out);
	reg32 r7428 (rst, clk, in, r7428_out);
	reg32 r7429 (rst, clk, in, r7429_out);
	reg32 r7430 (rst, clk, in, r7430_out);
	reg32 r7431 (rst, clk, in, r7431_out);
	reg32 r7432 (rst, clk, in, r7432_out);
	reg32 r7433 (rst, clk, in, r7433_out);
	reg32 r7434 (rst, clk, in, r7434_out);
	reg32 r7435 (rst, clk, in, r7435_out);
	reg32 r7436 (rst, clk, in, r7436_out);
	reg32 r7437 (rst, clk, in, r7437_out);
	reg32 r7438 (rst, clk, in, r7438_out);
	reg32 r7439 (rst, clk, in, r7439_out);
	reg32 r7440 (rst, clk, in, r7440_out);
	reg32 r7441 (rst, clk, in, r7441_out);
	reg32 r7442 (rst, clk, in, r7442_out);
	reg32 r7443 (rst, clk, in, r7443_out);
	reg32 r7444 (rst, clk, in, r7444_out);
	reg32 r7445 (rst, clk, in, r7445_out);
	reg32 r7446 (rst, clk, in, r7446_out);
	reg32 r7447 (rst, clk, in, r7447_out);
	reg32 r7448 (rst, clk, in, r7448_out);
	reg32 r7449 (rst, clk, in, r7449_out);
	reg32 r7450 (rst, clk, in, r7450_out);
	reg32 r7451 (rst, clk, in, r7451_out);
	reg32 r7452 (rst, clk, in, r7452_out);
	reg32 r7453 (rst, clk, in, r7453_out);
	reg32 r7454 (rst, clk, in, r7454_out);
	reg32 r7455 (rst, clk, in, r7455_out);
	reg32 r7456 (rst, clk, in, r7456_out);
	reg32 r7457 (rst, clk, in, r7457_out);
	reg32 r7458 (rst, clk, in, r7458_out);
	reg32 r7459 (rst, clk, in, r7459_out);
	reg32 r7460 (rst, clk, in, r7460_out);
	reg32 r7461 (rst, clk, in, r7461_out);
	reg32 r7462 (rst, clk, in, r7462_out);
	reg32 r7463 (rst, clk, in, r7463_out);
	reg32 r7464 (rst, clk, in, r7464_out);
	reg32 r7465 (rst, clk, in, r7465_out);
	reg32 r7466 (rst, clk, in, r7466_out);
	reg32 r7467 (rst, clk, in, r7467_out);
	reg32 r7468 (rst, clk, in, r7468_out);
	reg32 r7469 (rst, clk, in, r7469_out);
	reg32 r7470 (rst, clk, in, r7470_out);
	reg32 r7471 (rst, clk, in, r7471_out);
	reg32 r7472 (rst, clk, in, r7472_out);
	reg32 r7473 (rst, clk, in, r7473_out);
	reg32 r7474 (rst, clk, in, r7474_out);
	reg32 r7475 (rst, clk, in, r7475_out);
	reg32 r7476 (rst, clk, in, r7476_out);
	reg32 r7477 (rst, clk, in, r7477_out);
	reg32 r7478 (rst, clk, in, r7478_out);
	reg32 r7479 (rst, clk, in, r7479_out);
	reg32 r7480 (rst, clk, in, r7480_out);
	reg32 r7481 (rst, clk, in, r7481_out);
	reg32 r7482 (rst, clk, in, r7482_out);
	reg32 r7483 (rst, clk, in, r7483_out);
	reg32 r7484 (rst, clk, in, r7484_out);
	reg32 r7485 (rst, clk, in, r7485_out);
	reg32 r7486 (rst, clk, in, r7486_out);
	reg32 r7487 (rst, clk, in, r7487_out);
	reg32 r7488 (rst, clk, in, r7488_out);
	reg32 r7489 (rst, clk, in, r7489_out);
	reg32 r7490 (rst, clk, in, r7490_out);
	reg32 r7491 (rst, clk, in, r7491_out);
	reg32 r7492 (rst, clk, in, r7492_out);
	reg32 r7493 (rst, clk, in, r7493_out);
	reg32 r7494 (rst, clk, in, r7494_out);
	reg32 r7495 (rst, clk, in, r7495_out);
	reg32 r7496 (rst, clk, in, r7496_out);
	reg32 r7497 (rst, clk, in, r7497_out);
	reg32 r7498 (rst, clk, in, r7498_out);
	reg32 r7499 (rst, clk, in, r7499_out);
	reg32 r7500 (rst, clk, in, r7500_out);
	reg32 r7501 (rst, clk, in, r7501_out);
	reg32 r7502 (rst, clk, in, r7502_out);
	reg32 r7503 (rst, clk, in, r7503_out);
	reg32 r7504 (rst, clk, in, r7504_out);
	reg32 r7505 (rst, clk, in, r7505_out);
	reg32 r7506 (rst, clk, in, r7506_out);
	reg32 r7507 (rst, clk, in, r7507_out);
	reg32 r7508 (rst, clk, in, r7508_out);
	reg32 r7509 (rst, clk, in, r7509_out);
	reg32 r7510 (rst, clk, in, r7510_out);
	reg32 r7511 (rst, clk, in, r7511_out);
	reg32 r7512 (rst, clk, in, r7512_out);
	reg32 r7513 (rst, clk, in, r7513_out);
	reg32 r7514 (rst, clk, in, r7514_out);
	reg32 r7515 (rst, clk, in, r7515_out);
	reg32 r7516 (rst, clk, in, r7516_out);
	reg32 r7517 (rst, clk, in, r7517_out);
	reg32 r7518 (rst, clk, in, r7518_out);
	reg32 r7519 (rst, clk, in, r7519_out);
	reg32 r7520 (rst, clk, in, r7520_out);
	reg32 r7521 (rst, clk, in, r7521_out);
	reg32 r7522 (rst, clk, in, r7522_out);
	reg32 r7523 (rst, clk, in, r7523_out);
	reg32 r7524 (rst, clk, in, r7524_out);
	reg32 r7525 (rst, clk, in, r7525_out);
	reg32 r7526 (rst, clk, in, r7526_out);
	reg32 r7527 (rst, clk, in, r7527_out);
	reg32 r7528 (rst, clk, in, r7528_out);
	reg32 r7529 (rst, clk, in, r7529_out);
	reg32 r7530 (rst, clk, in, r7530_out);
	reg32 r7531 (rst, clk, in, r7531_out);
	reg32 r7532 (rst, clk, in, r7532_out);
	reg32 r7533 (rst, clk, in, r7533_out);
	reg32 r7534 (rst, clk, in, r7534_out);
	reg32 r7535 (rst, clk, in, r7535_out);
	reg32 r7536 (rst, clk, in, r7536_out);
	reg32 r7537 (rst, clk, in, r7537_out);
	reg32 r7538 (rst, clk, in, r7538_out);
	reg32 r7539 (rst, clk, in, r7539_out);
	reg32 r7540 (rst, clk, in, r7540_out);
	reg32 r7541 (rst, clk, in, r7541_out);
	reg32 r7542 (rst, clk, in, r7542_out);
	reg32 r7543 (rst, clk, in, r7543_out);
	reg32 r7544 (rst, clk, in, r7544_out);
	reg32 r7545 (rst, clk, in, r7545_out);
	reg32 r7546 (rst, clk, in, r7546_out);
	reg32 r7547 (rst, clk, in, r7547_out);
	reg32 r7548 (rst, clk, in, r7548_out);
	reg32 r7549 (rst, clk, in, r7549_out);
	reg32 r7550 (rst, clk, in, r7550_out);
	reg32 r7551 (rst, clk, in, r7551_out);
	reg32 r7552 (rst, clk, in, r7552_out);
	reg32 r7553 (rst, clk, in, r7553_out);
	reg32 r7554 (rst, clk, in, r7554_out);
	reg32 r7555 (rst, clk, in, r7555_out);
	reg32 r7556 (rst, clk, in, r7556_out);
	reg32 r7557 (rst, clk, in, r7557_out);
	reg32 r7558 (rst, clk, in, r7558_out);
	reg32 r7559 (rst, clk, in, r7559_out);
	reg32 r7560 (rst, clk, in, r7560_out);
	reg32 r7561 (rst, clk, in, r7561_out);
	reg32 r7562 (rst, clk, in, r7562_out);
	reg32 r7563 (rst, clk, in, r7563_out);
	reg32 r7564 (rst, clk, in, r7564_out);
	reg32 r7565 (rst, clk, in, r7565_out);
	reg32 r7566 (rst, clk, in, r7566_out);
	reg32 r7567 (rst, clk, in, r7567_out);
	reg32 r7568 (rst, clk, in, r7568_out);
	reg32 r7569 (rst, clk, in, r7569_out);
	reg32 r7570 (rst, clk, in, r7570_out);
	reg32 r7571 (rst, clk, in, r7571_out);
	reg32 r7572 (rst, clk, in, r7572_out);
	reg32 r7573 (rst, clk, in, r7573_out);
	reg32 r7574 (rst, clk, in, r7574_out);
	reg32 r7575 (rst, clk, in, r7575_out);
	reg32 r7576 (rst, clk, in, r7576_out);
	reg32 r7577 (rst, clk, in, r7577_out);
	reg32 r7578 (rst, clk, in, r7578_out);
	reg32 r7579 (rst, clk, in, r7579_out);
	reg32 r7580 (rst, clk, in, r7580_out);
	reg32 r7581 (rst, clk, in, r7581_out);
	reg32 r7582 (rst, clk, in, r7582_out);
	reg32 r7583 (rst, clk, in, r7583_out);
	reg32 r7584 (rst, clk, in, r7584_out);
	reg32 r7585 (rst, clk, in, r7585_out);
	reg32 r7586 (rst, clk, in, r7586_out);
	reg32 r7587 (rst, clk, in, r7587_out);
	reg32 r7588 (rst, clk, in, r7588_out);
	reg32 r7589 (rst, clk, in, r7589_out);
	reg32 r7590 (rst, clk, in, r7590_out);
	reg32 r7591 (rst, clk, in, r7591_out);
	reg32 r7592 (rst, clk, in, r7592_out);
	reg32 r7593 (rst, clk, in, r7593_out);
	reg32 r7594 (rst, clk, in, r7594_out);
	reg32 r7595 (rst, clk, in, r7595_out);
	reg32 r7596 (rst, clk, in, r7596_out);
	reg32 r7597 (rst, clk, in, r7597_out);
	reg32 r7598 (rst, clk, in, r7598_out);
	reg32 r7599 (rst, clk, in, r7599_out);
	reg32 r7600 (rst, clk, in, r7600_out);
	reg32 r7601 (rst, clk, in, r7601_out);
	reg32 r7602 (rst, clk, in, r7602_out);
	reg32 r7603 (rst, clk, in, r7603_out);
	reg32 r7604 (rst, clk, in, r7604_out);
	reg32 r7605 (rst, clk, in, r7605_out);
	reg32 r7606 (rst, clk, in, r7606_out);
	reg32 r7607 (rst, clk, in, r7607_out);
	reg32 r7608 (rst, clk, in, r7608_out);
	reg32 r7609 (rst, clk, in, r7609_out);
	reg32 r7610 (rst, clk, in, r7610_out);
	reg32 r7611 (rst, clk, in, r7611_out);
	reg32 r7612 (rst, clk, in, r7612_out);
	reg32 r7613 (rst, clk, in, r7613_out);
	reg32 r7614 (rst, clk, in, r7614_out);
	reg32 r7615 (rst, clk, in, r7615_out);
	reg32 r7616 (rst, clk, in, r7616_out);
	reg32 r7617 (rst, clk, in, r7617_out);
	reg32 r7618 (rst, clk, in, r7618_out);
	reg32 r7619 (rst, clk, in, r7619_out);
	reg32 r7620 (rst, clk, in, r7620_out);
	reg32 r7621 (rst, clk, in, r7621_out);
	reg32 r7622 (rst, clk, in, r7622_out);
	reg32 r7623 (rst, clk, in, r7623_out);
	reg32 r7624 (rst, clk, in, r7624_out);
	reg32 r7625 (rst, clk, in, r7625_out);
	reg32 r7626 (rst, clk, in, r7626_out);
	reg32 r7627 (rst, clk, in, r7627_out);
	reg32 r7628 (rst, clk, in, r7628_out);
	reg32 r7629 (rst, clk, in, r7629_out);
	reg32 r7630 (rst, clk, in, r7630_out);
	reg32 r7631 (rst, clk, in, r7631_out);
	reg32 r7632 (rst, clk, in, r7632_out);
	reg32 r7633 (rst, clk, in, r7633_out);
	reg32 r7634 (rst, clk, in, r7634_out);
	reg32 r7635 (rst, clk, in, r7635_out);
	reg32 r7636 (rst, clk, in, r7636_out);
	reg32 r7637 (rst, clk, in, r7637_out);
	reg32 r7638 (rst, clk, in, r7638_out);
	reg32 r7639 (rst, clk, in, r7639_out);
	reg32 r7640 (rst, clk, in, r7640_out);
	reg32 r7641 (rst, clk, in, r7641_out);
	reg32 r7642 (rst, clk, in, r7642_out);
	reg32 r7643 (rst, clk, in, r7643_out);
	reg32 r7644 (rst, clk, in, r7644_out);
	reg32 r7645 (rst, clk, in, r7645_out);
	reg32 r7646 (rst, clk, in, r7646_out);
	reg32 r7647 (rst, clk, in, r7647_out);
	reg32 r7648 (rst, clk, in, r7648_out);
	reg32 r7649 (rst, clk, in, r7649_out);
	reg32 r7650 (rst, clk, in, r7650_out);
	reg32 r7651 (rst, clk, in, r7651_out);
	reg32 r7652 (rst, clk, in, r7652_out);
	reg32 r7653 (rst, clk, in, r7653_out);
	reg32 r7654 (rst, clk, in, r7654_out);
	reg32 r7655 (rst, clk, in, r7655_out);
	reg32 r7656 (rst, clk, in, r7656_out);
	reg32 r7657 (rst, clk, in, r7657_out);
	reg32 r7658 (rst, clk, in, r7658_out);
	reg32 r7659 (rst, clk, in, r7659_out);
	reg32 r7660 (rst, clk, in, r7660_out);
	reg32 r7661 (rst, clk, in, r7661_out);
	reg32 r7662 (rst, clk, in, r7662_out);
	reg32 r7663 (rst, clk, in, r7663_out);
	reg32 r7664 (rst, clk, in, r7664_out);
	reg32 r7665 (rst, clk, in, r7665_out);
	reg32 r7666 (rst, clk, in, r7666_out);
	reg32 r7667 (rst, clk, in, r7667_out);
	reg32 r7668 (rst, clk, in, r7668_out);
	reg32 r7669 (rst, clk, in, r7669_out);
	reg32 r7670 (rst, clk, in, r7670_out);
	reg32 r7671 (rst, clk, in, r7671_out);
	reg32 r7672 (rst, clk, in, r7672_out);
	reg32 r7673 (rst, clk, in, r7673_out);
	reg32 r7674 (rst, clk, in, r7674_out);
	reg32 r7675 (rst, clk, in, r7675_out);
	reg32 r7676 (rst, clk, in, r7676_out);
	reg32 r7677 (rst, clk, in, r7677_out);
	reg32 r7678 (rst, clk, in, r7678_out);
	reg32 r7679 (rst, clk, in, r7679_out);
	reg32 r7680 (rst, clk, in, r7680_out);
	reg32 r7681 (rst, clk, in, r7681_out);
	reg32 r7682 (rst, clk, in, r7682_out);
	reg32 r7683 (rst, clk, in, r7683_out);
	reg32 r7684 (rst, clk, in, r7684_out);
	reg32 r7685 (rst, clk, in, r7685_out);
	reg32 r7686 (rst, clk, in, r7686_out);
	reg32 r7687 (rst, clk, in, r7687_out);
	reg32 r7688 (rst, clk, in, r7688_out);
	reg32 r7689 (rst, clk, in, r7689_out);
	reg32 r7690 (rst, clk, in, r7690_out);
	reg32 r7691 (rst, clk, in, r7691_out);
	reg32 r7692 (rst, clk, in, r7692_out);
	reg32 r7693 (rst, clk, in, r7693_out);
	reg32 r7694 (rst, clk, in, r7694_out);
	reg32 r7695 (rst, clk, in, r7695_out);
	reg32 r7696 (rst, clk, in, r7696_out);
	reg32 r7697 (rst, clk, in, r7697_out);
	reg32 r7698 (rst, clk, in, r7698_out);
	reg32 r7699 (rst, clk, in, r7699_out);
	reg32 r7700 (rst, clk, in, r7700_out);
	reg32 r7701 (rst, clk, in, r7701_out);
	reg32 r7702 (rst, clk, in, r7702_out);
	reg32 r7703 (rst, clk, in, r7703_out);
	reg32 r7704 (rst, clk, in, r7704_out);
	reg32 r7705 (rst, clk, in, r7705_out);
	reg32 r7706 (rst, clk, in, r7706_out);
	reg32 r7707 (rst, clk, in, r7707_out);
	reg32 r7708 (rst, clk, in, r7708_out);
	reg32 r7709 (rst, clk, in, r7709_out);
	reg32 r7710 (rst, clk, in, r7710_out);
	reg32 r7711 (rst, clk, in, r7711_out);
	reg32 r7712 (rst, clk, in, r7712_out);
	reg32 r7713 (rst, clk, in, r7713_out);
	reg32 r7714 (rst, clk, in, r7714_out);
	reg32 r7715 (rst, clk, in, r7715_out);
	reg32 r7716 (rst, clk, in, r7716_out);
	reg32 r7717 (rst, clk, in, r7717_out);
	reg32 r7718 (rst, clk, in, r7718_out);
	reg32 r7719 (rst, clk, in, r7719_out);
	reg32 r7720 (rst, clk, in, r7720_out);
	reg32 r7721 (rst, clk, in, r7721_out);
	reg32 r7722 (rst, clk, in, r7722_out);
	reg32 r7723 (rst, clk, in, r7723_out);
	reg32 r7724 (rst, clk, in, r7724_out);
	reg32 r7725 (rst, clk, in, r7725_out);
	reg32 r7726 (rst, clk, in, r7726_out);
	reg32 r7727 (rst, clk, in, r7727_out);
	reg32 r7728 (rst, clk, in, r7728_out);
	reg32 r7729 (rst, clk, in, r7729_out);
	reg32 r7730 (rst, clk, in, r7730_out);
	reg32 r7731 (rst, clk, in, r7731_out);
	reg32 r7732 (rst, clk, in, r7732_out);
	reg32 r7733 (rst, clk, in, r7733_out);
	reg32 r7734 (rst, clk, in, r7734_out);
	reg32 r7735 (rst, clk, in, r7735_out);
	reg32 r7736 (rst, clk, in, r7736_out);
	reg32 r7737 (rst, clk, in, r7737_out);
	reg32 r7738 (rst, clk, in, r7738_out);
	reg32 r7739 (rst, clk, in, r7739_out);
	reg32 r7740 (rst, clk, in, r7740_out);
	reg32 r7741 (rst, clk, in, r7741_out);
	reg32 r7742 (rst, clk, in, r7742_out);
	reg32 r7743 (rst, clk, in, r7743_out);
	reg32 r7744 (rst, clk, in, r7744_out);
	reg32 r7745 (rst, clk, in, r7745_out);
	reg32 r7746 (rst, clk, in, r7746_out);
	reg32 r7747 (rst, clk, in, r7747_out);
	reg32 r7748 (rst, clk, in, r7748_out);
	reg32 r7749 (rst, clk, in, r7749_out);
	reg32 r7750 (rst, clk, in, r7750_out);
	reg32 r7751 (rst, clk, in, r7751_out);
	reg32 r7752 (rst, clk, in, r7752_out);
	reg32 r7753 (rst, clk, in, r7753_out);
	reg32 r7754 (rst, clk, in, r7754_out);
	reg32 r7755 (rst, clk, in, r7755_out);
	reg32 r7756 (rst, clk, in, r7756_out);
	reg32 r7757 (rst, clk, in, r7757_out);
	reg32 r7758 (rst, clk, in, r7758_out);
	reg32 r7759 (rst, clk, in, r7759_out);
	reg32 r7760 (rst, clk, in, r7760_out);
	reg32 r7761 (rst, clk, in, r7761_out);
	reg32 r7762 (rst, clk, in, r7762_out);
	reg32 r7763 (rst, clk, in, r7763_out);
	reg32 r7764 (rst, clk, in, r7764_out);
	reg32 r7765 (rst, clk, in, r7765_out);
	reg32 r7766 (rst, clk, in, r7766_out);
	reg32 r7767 (rst, clk, in, r7767_out);
	reg32 r7768 (rst, clk, in, r7768_out);
	reg32 r7769 (rst, clk, in, r7769_out);
	reg32 r7770 (rst, clk, in, r7770_out);
	reg32 r7771 (rst, clk, in, r7771_out);
	reg32 r7772 (rst, clk, in, r7772_out);
	reg32 r7773 (rst, clk, in, r7773_out);
	reg32 r7774 (rst, clk, in, r7774_out);
	reg32 r7775 (rst, clk, in, r7775_out);
	reg32 r7776 (rst, clk, in, r7776_out);
	reg32 r7777 (rst, clk, in, r7777_out);
	reg32 r7778 (rst, clk, in, r7778_out);
	reg32 r7779 (rst, clk, in, r7779_out);
	reg32 r7780 (rst, clk, in, r7780_out);
	reg32 r7781 (rst, clk, in, r7781_out);
	reg32 r7782 (rst, clk, in, r7782_out);
	reg32 r7783 (rst, clk, in, r7783_out);
	reg32 r7784 (rst, clk, in, r7784_out);
	reg32 r7785 (rst, clk, in, r7785_out);
	reg32 r7786 (rst, clk, in, r7786_out);
	reg32 r7787 (rst, clk, in, r7787_out);
	reg32 r7788 (rst, clk, in, r7788_out);
	reg32 r7789 (rst, clk, in, r7789_out);
	reg32 r7790 (rst, clk, in, r7790_out);
	reg32 r7791 (rst, clk, in, r7791_out);
	reg32 r7792 (rst, clk, in, r7792_out);
	reg32 r7793 (rst, clk, in, r7793_out);
	reg32 r7794 (rst, clk, in, r7794_out);
	reg32 r7795 (rst, clk, in, r7795_out);
	reg32 r7796 (rst, clk, in, r7796_out);
	reg32 r7797 (rst, clk, in, r7797_out);
	reg32 r7798 (rst, clk, in, r7798_out);
	reg32 r7799 (rst, clk, in, r7799_out);
	reg32 r7800 (rst, clk, in, r7800_out);
	reg32 r7801 (rst, clk, in, r7801_out);
	reg32 r7802 (rst, clk, in, r7802_out);
	reg32 r7803 (rst, clk, in, r7803_out);
	reg32 r7804 (rst, clk, in, r7804_out);
	reg32 r7805 (rst, clk, in, r7805_out);
	reg32 r7806 (rst, clk, in, r7806_out);
	reg32 r7807 (rst, clk, in, r7807_out);
	reg32 r7808 (rst, clk, in, r7808_out);
	reg32 r7809 (rst, clk, in, r7809_out);
	reg32 r7810 (rst, clk, in, r7810_out);
	reg32 r7811 (rst, clk, in, r7811_out);
	reg32 r7812 (rst, clk, in, r7812_out);
	reg32 r7813 (rst, clk, in, r7813_out);
	reg32 r7814 (rst, clk, in, r7814_out);
	reg32 r7815 (rst, clk, in, r7815_out);
	reg32 r7816 (rst, clk, in, r7816_out);
	reg32 r7817 (rst, clk, in, r7817_out);
	reg32 r7818 (rst, clk, in, r7818_out);
	reg32 r7819 (rst, clk, in, r7819_out);
	reg32 r7820 (rst, clk, in, r7820_out);
	reg32 r7821 (rst, clk, in, r7821_out);
	reg32 r7822 (rst, clk, in, r7822_out);
	reg32 r7823 (rst, clk, in, r7823_out);
	reg32 r7824 (rst, clk, in, r7824_out);
	reg32 r7825 (rst, clk, in, r7825_out);
	reg32 r7826 (rst, clk, in, r7826_out);
	reg32 r7827 (rst, clk, in, r7827_out);
	reg32 r7828 (rst, clk, in, r7828_out);
	reg32 r7829 (rst, clk, in, r7829_out);
	reg32 r7830 (rst, clk, in, r7830_out);
	reg32 r7831 (rst, clk, in, r7831_out);
	reg32 r7832 (rst, clk, in, r7832_out);
	reg32 r7833 (rst, clk, in, r7833_out);
	reg32 r7834 (rst, clk, in, r7834_out);
	reg32 r7835 (rst, clk, in, r7835_out);
	reg32 r7836 (rst, clk, in, r7836_out);
	reg32 r7837 (rst, clk, in, r7837_out);
	reg32 r7838 (rst, clk, in, r7838_out);
	reg32 r7839 (rst, clk, in, r7839_out);
	reg32 r7840 (rst, clk, in, r7840_out);
	reg32 r7841 (rst, clk, in, r7841_out);
	reg32 r7842 (rst, clk, in, r7842_out);
	reg32 r7843 (rst, clk, in, r7843_out);
	reg32 r7844 (rst, clk, in, r7844_out);
	reg32 r7845 (rst, clk, in, r7845_out);
	reg32 r7846 (rst, clk, in, r7846_out);
	reg32 r7847 (rst, clk, in, r7847_out);
	reg32 r7848 (rst, clk, in, r7848_out);
	reg32 r7849 (rst, clk, in, r7849_out);
	reg32 r7850 (rst, clk, in, r7850_out);
	reg32 r7851 (rst, clk, in, r7851_out);
	reg32 r7852 (rst, clk, in, r7852_out);
	reg32 r7853 (rst, clk, in, r7853_out);
	reg32 r7854 (rst, clk, in, r7854_out);
	reg32 r7855 (rst, clk, in, r7855_out);
	reg32 r7856 (rst, clk, in, r7856_out);
	reg32 r7857 (rst, clk, in, r7857_out);
	reg32 r7858 (rst, clk, in, r7858_out);
	reg32 r7859 (rst, clk, in, r7859_out);
	reg32 r7860 (rst, clk, in, r7860_out);
	reg32 r7861 (rst, clk, in, r7861_out);
	reg32 r7862 (rst, clk, in, r7862_out);
	reg32 r7863 (rst, clk, in, r7863_out);
	reg32 r7864 (rst, clk, in, r7864_out);
	reg32 r7865 (rst, clk, in, r7865_out);
	reg32 r7866 (rst, clk, in, r7866_out);
	reg32 r7867 (rst, clk, in, r7867_out);
	reg32 r7868 (rst, clk, in, r7868_out);
	reg32 r7869 (rst, clk, in, r7869_out);
	reg32 r7870 (rst, clk, in, r7870_out);
	reg32 r7871 (rst, clk, in, r7871_out);
	reg32 r7872 (rst, clk, in, r7872_out);
	reg32 r7873 (rst, clk, in, r7873_out);
	reg32 r7874 (rst, clk, in, r7874_out);
	reg32 r7875 (rst, clk, in, r7875_out);
	reg32 r7876 (rst, clk, in, r7876_out);
	reg32 r7877 (rst, clk, in, r7877_out);
	reg32 r7878 (rst, clk, in, r7878_out);
	reg32 r7879 (rst, clk, in, r7879_out);
	reg32 r7880 (rst, clk, in, r7880_out);
	reg32 r7881 (rst, clk, in, r7881_out);
	reg32 r7882 (rst, clk, in, r7882_out);
	reg32 r7883 (rst, clk, in, r7883_out);
	reg32 r7884 (rst, clk, in, r7884_out);
	reg32 r7885 (rst, clk, in, r7885_out);
	reg32 r7886 (rst, clk, in, r7886_out);
	reg32 r7887 (rst, clk, in, r7887_out);
	reg32 r7888 (rst, clk, in, r7888_out);
	reg32 r7889 (rst, clk, in, r7889_out);
	reg32 r7890 (rst, clk, in, r7890_out);
	reg32 r7891 (rst, clk, in, r7891_out);
	reg32 r7892 (rst, clk, in, r7892_out);
	reg32 r7893 (rst, clk, in, r7893_out);
	reg32 r7894 (rst, clk, in, r7894_out);
	reg32 r7895 (rst, clk, in, r7895_out);
	reg32 r7896 (rst, clk, in, r7896_out);
	reg32 r7897 (rst, clk, in, r7897_out);
	reg32 r7898 (rst, clk, in, r7898_out);
	reg32 r7899 (rst, clk, in, r7899_out);
	reg32 r7900 (rst, clk, in, r7900_out);
	reg32 r7901 (rst, clk, in, r7901_out);
	reg32 r7902 (rst, clk, in, r7902_out);
	reg32 r7903 (rst, clk, in, r7903_out);
	reg32 r7904 (rst, clk, in, r7904_out);
	reg32 r7905 (rst, clk, in, r7905_out);
	reg32 r7906 (rst, clk, in, r7906_out);
	reg32 r7907 (rst, clk, in, r7907_out);
	reg32 r7908 (rst, clk, in, r7908_out);
	reg32 r7909 (rst, clk, in, r7909_out);
	reg32 r7910 (rst, clk, in, r7910_out);
	reg32 r7911 (rst, clk, in, r7911_out);
	reg32 r7912 (rst, clk, in, r7912_out);
	reg32 r7913 (rst, clk, in, r7913_out);
	reg32 r7914 (rst, clk, in, r7914_out);
	reg32 r7915 (rst, clk, in, r7915_out);
	reg32 r7916 (rst, clk, in, r7916_out);
	reg32 r7917 (rst, clk, in, r7917_out);
	reg32 r7918 (rst, clk, in, r7918_out);
	reg32 r7919 (rst, clk, in, r7919_out);
	reg32 r7920 (rst, clk, in, r7920_out);
	reg32 r7921 (rst, clk, in, r7921_out);
	reg32 r7922 (rst, clk, in, r7922_out);
	reg32 r7923 (rst, clk, in, r7923_out);
	reg32 r7924 (rst, clk, in, r7924_out);
	reg32 r7925 (rst, clk, in, r7925_out);
	reg32 r7926 (rst, clk, in, r7926_out);
	reg32 r7927 (rst, clk, in, r7927_out);
	reg32 r7928 (rst, clk, in, r7928_out);
	reg32 r7929 (rst, clk, in, r7929_out);
	reg32 r7930 (rst, clk, in, r7930_out);
	reg32 r7931 (rst, clk, in, r7931_out);
	reg32 r7932 (rst, clk, in, r7932_out);
	reg32 r7933 (rst, clk, in, r7933_out);
	reg32 r7934 (rst, clk, in, r7934_out);
	reg32 r7935 (rst, clk, in, r7935_out);
	reg32 r7936 (rst, clk, in, r7936_out);
	reg32 r7937 (rst, clk, in, r7937_out);
	reg32 r7938 (rst, clk, in, r7938_out);
	reg32 r7939 (rst, clk, in, r7939_out);
	reg32 r7940 (rst, clk, in, r7940_out);
	reg32 r7941 (rst, clk, in, r7941_out);
	reg32 r7942 (rst, clk, in, r7942_out);
	reg32 r7943 (rst, clk, in, r7943_out);
	reg32 r7944 (rst, clk, in, r7944_out);
	reg32 r7945 (rst, clk, in, r7945_out);
	reg32 r7946 (rst, clk, in, r7946_out);
	reg32 r7947 (rst, clk, in, r7947_out);
	reg32 r7948 (rst, clk, in, r7948_out);
	reg32 r7949 (rst, clk, in, r7949_out);
	reg32 r7950 (rst, clk, in, r7950_out);
	reg32 r7951 (rst, clk, in, r7951_out);
	reg32 r7952 (rst, clk, in, r7952_out);
	reg32 r7953 (rst, clk, in, r7953_out);
	reg32 r7954 (rst, clk, in, r7954_out);
	reg32 r7955 (rst, clk, in, r7955_out);
	reg32 r7956 (rst, clk, in, r7956_out);
	reg32 r7957 (rst, clk, in, r7957_out);
	reg32 r7958 (rst, clk, in, r7958_out);
	reg32 r7959 (rst, clk, in, r7959_out);
	reg32 r7960 (rst, clk, in, r7960_out);
	reg32 r7961 (rst, clk, in, r7961_out);
	reg32 r7962 (rst, clk, in, r7962_out);
	reg32 r7963 (rst, clk, in, r7963_out);
	reg32 r7964 (rst, clk, in, r7964_out);
	reg32 r7965 (rst, clk, in, r7965_out);
	reg32 r7966 (rst, clk, in, r7966_out);
	reg32 r7967 (rst, clk, in, r7967_out);
	reg32 r7968 (rst, clk, in, r7968_out);
	reg32 r7969 (rst, clk, in, r7969_out);
	reg32 r7970 (rst, clk, in, r7970_out);
	reg32 r7971 (rst, clk, in, r7971_out);
	reg32 r7972 (rst, clk, in, r7972_out);
	reg32 r7973 (rst, clk, in, r7973_out);
	reg32 r7974 (rst, clk, in, r7974_out);
	reg32 r7975 (rst, clk, in, r7975_out);
	reg32 r7976 (rst, clk, in, r7976_out);
	reg32 r7977 (rst, clk, in, r7977_out);
	reg32 r7978 (rst, clk, in, r7978_out);
	reg32 r7979 (rst, clk, in, r7979_out);
	reg32 r7980 (rst, clk, in, r7980_out);
	reg32 r7981 (rst, clk, in, r7981_out);
	reg32 r7982 (rst, clk, in, r7982_out);
	reg32 r7983 (rst, clk, in, r7983_out);
	reg32 r7984 (rst, clk, in, r7984_out);
	reg32 r7985 (rst, clk, in, r7985_out);
	reg32 r7986 (rst, clk, in, r7986_out);
	reg32 r7987 (rst, clk, in, r7987_out);
	reg32 r7988 (rst, clk, in, r7988_out);
	reg32 r7989 (rst, clk, in, r7989_out);
	reg32 r7990 (rst, clk, in, r7990_out);
	reg32 r7991 (rst, clk, in, r7991_out);
	reg32 r7992 (rst, clk, in, r7992_out);
	reg32 r7993 (rst, clk, in, r7993_out);
	reg32 r7994 (rst, clk, in, r7994_out);
	reg32 r7995 (rst, clk, in, r7995_out);
	reg32 r7996 (rst, clk, in, r7996_out);
	reg32 r7997 (rst, clk, in, r7997_out);
	reg32 r7998 (rst, clk, in, r7998_out);
	reg32 r7999 (rst, clk, in, r7999_out);

	assign out = r7999_out;
endmodule
