-- Syndrome Error Correction Module.
--
-- This module attempts to apply Syndrome error correction to the input
-- encoded vector.
-- This module effectively assumes we have received our received_codeword
-- which has possible errors in it. It calculates the syndrome of the
-- codeword and applies the syndrome (assuming we find one that is in our
-- known set) to the codeword. Finaly it extracts the message. 
--
-- Author: Malcolm Watt

library ieee;
use ieee.std_logic_1164.all;


entity syndrome_correction is
	port(
		received_codeword : in std_logic_vector(15 downto 0);
		decoded_message : out std_logic_vector(4 downto 0)
	);
end syndrome_correction;


architecture corr of syndrome_correction is
	type H_matrix is array(15 downto 0, 10 downto 0) of std_logic;
	signal syndrome : std_logic_vector(10 downto 0) := (others => '0');
	signal error_vector : std_logic_vector(15 downto 0) := (others => '0');
	signal decoded_codeword : std_logic_vector(15 downto 0) := (others => '0');
	signal H_transpose : H_matrix;
	
	-- Hardcoded constant for the H matrix. This is actually the transpose of H.
	constant H_matrix_init : H_matrix:= (
		('1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '1'),
		('1', '1', '1', '0', '0', '0', '1', '1', '1', '0', '1'),
		('1', '0', '0', '1', '1', '0', '1', '1', '0', '1', '1'),
		('0', '1', '0', '1', '0', '1', '1', '0', '1', '1', '1'),
		('0', '0', '1', '0', '1', '1', '0', '1', '1', '1', '1'),
		('1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0'),
		('0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0'),
		('0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0'),
		('0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0'),
		('0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0'),
		('0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0'),
		('0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0'),
		('0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0'),
		('0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0'),
		('0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0'),
		('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1')
	);

	-- Get the syndrome. This function basically performs vector * matrix
	-- multiplication. Effectively the formula is synd = code_arg * H_arg
	-- which when we look back at our matlab implementation, is equivalent
	-- to our `syndrome = r * H';` line.
	function get_synd(H_arg : H_matrix; code_arg : std_logic_vector(15 downto 0))
	return std_logic_vector is
		variable synd : std_logic_vector(10 downto 0) := (others => '0');
	begin
		
		-- For each of the results, we XOR the result of ANDing the entries of the
		-- code_arg with the current columns values.
		for i in synd'range loop
			for j in 0 to 15 loop
				synd(i) := synd(i) XOR (code_arg(j) AND H_arg(j, i));
			end loop;
		end loop;
		return synd;
	end get_synd;

begin	
	H_transpose <= H_matrix_init; -- Set the H matrix (it is a constant array).
	
	-- Get the syndrome for the received_codeword and the H matrix.
	syndrome <= get_synd(H_transpose, received_codeword);
	
	-- Get the decoded_message by XORing and taking the first 5 bits.
	decoded_codeword <= received_codeword XOR error_vector;
	decoded_message <= decoded_codeword(4 downto 0);
	
	
	-- Figure out what the error_vector is based on the syndrome table.
	-- This is purely combinational logic. The cases were automatically
	-- generated by the print_syndrome_pairs matlab script found in
	-- the matlab directory.
	P1 : process(received_codeword, decoded_codeword) is
	begin
		check_syndromes : case syndrome is
			when "00000000000" => error_vector <= "0000000000000000";
			when "11111100001" => error_vector <= "1000000000000000";
			when "11100011101" => error_vector <= "0100000000000000";
			when "10011011011" => error_vector <= "0010000000000000";
			when "01010110111" => error_vector <= "0001000000000000";
			when "00101101111" => error_vector <= "0000100000000000";
			when "10000000000" => error_vector <= "0000010000000000";
			when "01000000000" => error_vector <= "0000001000000000";
			when "00100000000" => error_vector <= "0000000100000000";
			when "00010000000" => error_vector <= "0000000010000000";
			when "00001000000" => error_vector <= "0000000001000000";
			when "00000100000" => error_vector <= "0000000000100000";
			when "00000010000" => error_vector <= "0000000000010000";
			when "00000001000" => error_vector <= "0000000000001000";
			when "00000000100" => error_vector <= "0000000000000100";
			when "00000000010" => error_vector <= "0000000000000010";
			when "00000000001" => error_vector <= "0000000000000001";
			when "00011111100" => error_vector <= "1100000000000000";
			when "01100111010" => error_vector <= "1010000000000000";
			when "10101010110" => error_vector <= "1001000000000000";
			when "11010001110" => error_vector <= "1000100000000000";
			when "01111100001" => error_vector <= "1000010000000000";
			when "10111100001" => error_vector <= "1000001000000000";
			when "11011100001" => error_vector <= "1000000100000000";
			when "11101100001" => error_vector <= "1000000010000000";
			when "11110100001" => error_vector <= "1000000001000000";
			when "11111000001" => error_vector <= "1000000000100000";
			when "11111110001" => error_vector <= "1000000000010000";
			when "11111101001" => error_vector <= "1000000000001000";
			when "11111100101" => error_vector <= "1000000000000100";
			when "11111100011" => error_vector <= "1000000000000010";
			when "11111100000" => error_vector <= "1000000000000001";
			when "01111000110" => error_vector <= "0110000000000000";
			when "10110101010" => error_vector <= "0101000000000000";
			when "11001110010" => error_vector <= "0100100000000000";
			when "01100011101" => error_vector <= "0100010000000000";
			when "10100011101" => error_vector <= "0100001000000000";
			when "11000011101" => error_vector <= "0100000100000000";
			when "11110011101" => error_vector <= "0100000010000000";
			when "11101011101" => error_vector <= "0100000001000000";
			when "11100111101" => error_vector <= "0100000000100000";
			when "11100001101" => error_vector <= "0100000000010000";
			when "11100010101" => error_vector <= "0100000000001000";
			when "11100011001" => error_vector <= "0100000000000100";
			when "11100011111" => error_vector <= "0100000000000010";
			when "11100011100" => error_vector <= "0100000000000001";
			when "11001101100" => error_vector <= "0011000000000000";
			when "10110110100" => error_vector <= "0010100000000000";
			when "00011011011" => error_vector <= "0010010000000000";
			when "11011011011" => error_vector <= "0010001000000000";
			when "10111011011" => error_vector <= "0010000100000000";
			when "10001011011" => error_vector <= "0010000010000000";
			when "10010011011" => error_vector <= "0010000001000000";
			when "10011111011" => error_vector <= "0010000000100000";
			when "10011001011" => error_vector <= "0010000000010000";
			when "10011010011" => error_vector <= "0010000000001000";
			when "10011011111" => error_vector <= "0010000000000100";
			when "10011011001" => error_vector <= "0010000000000010";
			when "10011011010" => error_vector <= "0010000000000001";
			when "01111011000" => error_vector <= "0001100000000000";
			when "11010110111" => error_vector <= "0001010000000000";
			when "00010110111" => error_vector <= "0001001000000000";
			when "01110110111" => error_vector <= "0001000100000000";
			when "01000110111" => error_vector <= "0001000010000000";
			when "01011110111" => error_vector <= "0001000001000000";
			when "01010010111" => error_vector <= "0001000000100000";
			when "01010100111" => error_vector <= "0001000000010000";
			when "01010111111" => error_vector <= "0001000000001000";
			when "01010110011" => error_vector <= "0001000000000100";
			when "01010110101" => error_vector <= "0001000000000010";
			when "01010110110" => error_vector <= "0001000000000001";
			when "10101101111" => error_vector <= "0000110000000000";
			when "01101101111" => error_vector <= "0000101000000000";
			when "00001101111" => error_vector <= "0000100100000000";
			when "00111101111" => error_vector <= "0000100010000000";
			when "00100101111" => error_vector <= "0000100001000000";
			when "00101001111" => error_vector <= "0000100000100000";
			when "00101111111" => error_vector <= "0000100000010000";
			when "00101100111" => error_vector <= "0000100000001000";
			when "00101101011" => error_vector <= "0000100000000100";
			when "00101101101" => error_vector <= "0000100000000010";
			when "00101101110" => error_vector <= "0000100000000001";
			when "11000000000" => error_vector <= "0000011000000000";
			when "10100000000" => error_vector <= "0000010100000000";
			when "10010000000" => error_vector <= "0000010010000000";
			when "10001000000" => error_vector <= "0000010001000000";
			when "10000100000" => error_vector <= "0000010000100000";
			when "10000010000" => error_vector <= "0000010000010000";
			when "10000001000" => error_vector <= "0000010000001000";
			when "10000000100" => error_vector <= "0000010000000100";
			when "10000000010" => error_vector <= "0000010000000010";
			when "10000000001" => error_vector <= "0000010000000001";
			when "01100000000" => error_vector <= "0000001100000000";
			when "01010000000" => error_vector <= "0000001010000000";
			when "01001000000" => error_vector <= "0000001001000000";
			when "01000100000" => error_vector <= "0000001000100000";
			when "01000010000" => error_vector <= "0000001000010000";
			when "01000001000" => error_vector <= "0000001000001000";
			when "01000000100" => error_vector <= "0000001000000100";
			when "01000000010" => error_vector <= "0000001000000010";
			when "01000000001" => error_vector <= "0000001000000001";
			when "00110000000" => error_vector <= "0000000110000000";
			when "00101000000" => error_vector <= "0000000101000000";
			when "00100100000" => error_vector <= "0000000100100000";
			when "00100010000" => error_vector <= "0000000100010000";
			when "00100001000" => error_vector <= "0000000100001000";
			when "00100000100" => error_vector <= "0000000100000100";
			when "00100000010" => error_vector <= "0000000100000010";
			when "00100000001" => error_vector <= "0000000100000001";
			when "00011000000" => error_vector <= "0000000011000000";
			when "00010100000" => error_vector <= "0000000010100000";
			when "00010010000" => error_vector <= "0000000010010000";
			when "00010001000" => error_vector <= "0000000010001000";
			when "00010000100" => error_vector <= "0000000010000100";
			when "00010000010" => error_vector <= "0000000010000010";
			when "00010000001" => error_vector <= "0000000010000001";
			when "00001100000" => error_vector <= "0000000001100000";
			when "00001010000" => error_vector <= "0000000001010000";
			when "00001001000" => error_vector <= "0000000001001000";
			when "00001000100" => error_vector <= "0000000001000100";
			when "00001000010" => error_vector <= "0000000001000010";
			when "00001000001" => error_vector <= "0000000001000001";
			when "00000110000" => error_vector <= "0000000000110000";
			when "00000101000" => error_vector <= "0000000000101000";
			when "00000100100" => error_vector <= "0000000000100100";
			when "00000100010" => error_vector <= "0000000000100010";
			when "00000100001" => error_vector <= "0000000000100001";
			when "00000011000" => error_vector <= "0000000000011000";
			when "00000010100" => error_vector <= "0000000000010100";
			when "00000010010" => error_vector <= "0000000000010010";
			when "00000010001" => error_vector <= "0000000000010001";
			when "00000001100" => error_vector <= "0000000000001100";
			when "00000001010" => error_vector <= "0000000000001010";
			when "00000001001" => error_vector <= "0000000000001001";
			when "00000000110" => error_vector <= "0000000000000110";
			when "00000000101" => error_vector <= "0000000000000101";
			when "00000000011" => error_vector <= "0000000000000011";
			when "10000100111" => error_vector <= "1110000000000000";
			when "01001001011" => error_vector <= "1101000000000000";
			when "00110010011" => error_vector <= "1100100000000000";
			when "10011111100" => error_vector <= "1100010000000000";
			when "01011111100" => error_vector <= "1100001000000000";
			when "00111111100" => error_vector <= "1100000100000000";
			when "00001111100" => error_vector <= "1100000010000000";
			when "00010111100" => error_vector <= "1100000001000000";
			when "00011011100" => error_vector <= "1100000000100000";
			when "00011101100" => error_vector <= "1100000000010000";
			when "00011110100" => error_vector <= "1100000000001000";
			when "00011111000" => error_vector <= "1100000000000100";
			when "00011111110" => error_vector <= "1100000000000010";
			when "00011111101" => error_vector <= "1100000000000001";
			when "00110001101" => error_vector <= "1011000000000000";
			when "01001010101" => error_vector <= "1010100000000000";
			when "11100111010" => error_vector <= "1010010000000000";
			when "00100111010" => error_vector <= "1010001000000000";
			when "01000111010" => error_vector <= "1010000100000000";
			when "01110111010" => error_vector <= "1010000010000000";
			when "01101111010" => error_vector <= "1010000001000000";
			when "01100011010" => error_vector <= "1010000000100000";
			when "01100101010" => error_vector <= "1010000000010000";
			when "01100110010" => error_vector <= "1010000000001000";
			when "01100111110" => error_vector <= "1010000000000100";
			when "01100111000" => error_vector <= "1010000000000010";
			when "01100111011" => error_vector <= "1010000000000001";
			when "10000111001" => error_vector <= "1001100000000000";
			when "00101010110" => error_vector <= "1001010000000000";
			when "11101010110" => error_vector <= "1001001000000000";
			when "10001010110" => error_vector <= "1001000100000000";
			when "10111010110" => error_vector <= "1001000010000000";
			when "10100010110" => error_vector <= "1001000001000000";
			when "10101110110" => error_vector <= "1001000000100000";
			when "10101000110" => error_vector <= "1001000000010000";
			when "10101011110" => error_vector <= "1001000000001000";
			when "10101010010" => error_vector <= "1001000000000100";
			when "10101010100" => error_vector <= "1001000000000010";
			when "10101010111" => error_vector <= "1001000000000001";
			when "01010001110" => error_vector <= "1000110000000000";
			when "10010001110" => error_vector <= "1000101000000000";
			when "11110001110" => error_vector <= "1000100100000000";
			when "11000001110" => error_vector <= "1000100010000000";
			when "11011001110" => error_vector <= "1000100001000000";
			when "11010101110" => error_vector <= "1000100000100000";
			when "11010011110" => error_vector <= "1000100000010000";
			when "11010000110" => error_vector <= "1000100000001000";
			when "11010001010" => error_vector <= "1000100000000100";
			when "11010001100" => error_vector <= "1000100000000010";
			when "11010001111" => error_vector <= "1000100000000001";
			when "00111100001" => error_vector <= "1000011000000000";
			when "01011100001" => error_vector <= "1000010100000000";
			when "01101100001" => error_vector <= "1000010010000000";
			when "01110100001" => error_vector <= "1000010001000000";
			when "01111000001" => error_vector <= "1000010000100000";
			when "01111110001" => error_vector <= "1000010000010000";
			when "01111101001" => error_vector <= "1000010000001000";
			when "01111100101" => error_vector <= "1000010000000100";
			when "01111100011" => error_vector <= "1000010000000010";
			when "01111100000" => error_vector <= "1000010000000001";
			when "10011100001" => error_vector <= "1000001100000000";
			when "10101100001" => error_vector <= "1000001010000000";
			when "10110100001" => error_vector <= "1000001001000000";
			when "10111000001" => error_vector <= "1000001000100000";
			when "10111110001" => error_vector <= "1000001000010000";
			when "10111101001" => error_vector <= "1000001000001000";
			when "10111100101" => error_vector <= "1000001000000100";
			when "10111100011" => error_vector <= "1000001000000010";
			when "10111100000" => error_vector <= "1000001000000001";
			when "11001100001" => error_vector <= "1000000110000000";
			when "11010100001" => error_vector <= "1000000101000000";
			when "11011000001" => error_vector <= "1000000100100000";
			when "11011110001" => error_vector <= "1000000100010000";
			when "11011101001" => error_vector <= "1000000100001000";
			when "11011100101" => error_vector <= "1000000100000100";
			when "11011100011" => error_vector <= "1000000100000010";
			when "11011100000" => error_vector <= "1000000100000001";
			when "11100100001" => error_vector <= "1000000011000000";
			when "11101000001" => error_vector <= "1000000010100000";
			when "11101110001" => error_vector <= "1000000010010000";
			when "11101101001" => error_vector <= "1000000010001000";
			when "11101100101" => error_vector <= "1000000010000100";
			when "11101100011" => error_vector <= "1000000010000010";
			when "11101100000" => error_vector <= "1000000010000001";
			when "11110000001" => error_vector <= "1000000001100000";
			when "11110110001" => error_vector <= "1000000001010000";
			when "11110101001" => error_vector <= "1000000001001000";
			when "11110100101" => error_vector <= "1000000001000100";
			when "11110100011" => error_vector <= "1000000001000010";
			when "11110100000" => error_vector <= "1000000001000001";
			when "11111010001" => error_vector <= "1000000000110000";
			when "11111001001" => error_vector <= "1000000000101000";
			when "11111000101" => error_vector <= "1000000000100100";
			when "11111000011" => error_vector <= "1000000000100010";
			when "11111000000" => error_vector <= "1000000000100001";
			when "11111111001" => error_vector <= "1000000000011000";
			when "11111110101" => error_vector <= "1000000000010100";
			when "11111110011" => error_vector <= "1000000000010010";
			when "11111110000" => error_vector <= "1000000000010001";
			when "11111101101" => error_vector <= "1000000000001100";
			when "11111101011" => error_vector <= "1000000000001010";
			when "11111101000" => error_vector <= "1000000000001001";
			when "11111100111" => error_vector <= "1000000000000110";
			when "11111100100" => error_vector <= "1000000000000101";
			when "11111100010" => error_vector <= "1000000000000011";
			when "00101110001" => error_vector <= "0111000000000000";
			when "01010101001" => error_vector <= "0110100000000000";
			when "11111000110" => error_vector <= "0110010000000000";
			when "00111000110" => error_vector <= "0110001000000000";
			when "01011000110" => error_vector <= "0110000100000000";
			when "01101000110" => error_vector <= "0110000010000000";
			when "01110000110" => error_vector <= "0110000001000000";
			when "01111100110" => error_vector <= "0110000000100000";
			when "01111010110" => error_vector <= "0110000000010000";
			when "01111001110" => error_vector <= "0110000000001000";
			when "01111000010" => error_vector <= "0110000000000100";
			when "01111000100" => error_vector <= "0110000000000010";
			when "01111000111" => error_vector <= "0110000000000001";
			when "10011000101" => error_vector <= "0101100000000000";
			when "00110101010" => error_vector <= "0101010000000000";
			when "11110101010" => error_vector <= "0101001000000000";
			when "10010101010" => error_vector <= "0101000100000000";
			when "10100101010" => error_vector <= "0101000010000000";
			when "10111101010" => error_vector <= "0101000001000000";
			when "10110001010" => error_vector <= "0101000000100000";
			when "10110111010" => error_vector <= "0101000000010000";
			when "10110100010" => error_vector <= "0101000000001000";
			when "10110101110" => error_vector <= "0101000000000100";
			when "10110101000" => error_vector <= "0101000000000010";
			when "10110101011" => error_vector <= "0101000000000001";
			when "01001110010" => error_vector <= "0100110000000000";
			when "10001110010" => error_vector <= "0100101000000000";
			when "11101110010" => error_vector <= "0100100100000000";
			when "11011110010" => error_vector <= "0100100010000000";
			when "11000110010" => error_vector <= "0100100001000000";
			when "11001010010" => error_vector <= "0100100000100000";
			when "11001100010" => error_vector <= "0100100000010000";
			when "11001111010" => error_vector <= "0100100000001000";
			when "11001110110" => error_vector <= "0100100000000100";
			when "11001110000" => error_vector <= "0100100000000010";
			when "11001110011" => error_vector <= "0100100000000001";
			when "00100011101" => error_vector <= "0100011000000000";
			when "01000011101" => error_vector <= "0100010100000000";
			when "01110011101" => error_vector <= "0100010010000000";
			when "01101011101" => error_vector <= "0100010001000000";
			when "01100111101" => error_vector <= "0100010000100000";
			when "01100001101" => error_vector <= "0100010000010000";
			when "01100010101" => error_vector <= "0100010000001000";
			when "01100011001" => error_vector <= "0100010000000100";
			when "01100011111" => error_vector <= "0100010000000010";
			when "01100011100" => error_vector <= "0100010000000001";
			when "10000011101" => error_vector <= "0100001100000000";
			when "10110011101" => error_vector <= "0100001010000000";
			when "10101011101" => error_vector <= "0100001001000000";
			when "10100111101" => error_vector <= "0100001000100000";
			when "10100001101" => error_vector <= "0100001000010000";
			when "10100010101" => error_vector <= "0100001000001000";
			when "10100011001" => error_vector <= "0100001000000100";
			when "10100011111" => error_vector <= "0100001000000010";
			when "10100011100" => error_vector <= "0100001000000001";
			when "11010011101" => error_vector <= "0100000110000000";
			when "11001011101" => error_vector <= "0100000101000000";
			when "11000111101" => error_vector <= "0100000100100000";
			when "11000001101" => error_vector <= "0100000100010000";
			when "11000010101" => error_vector <= "0100000100001000";
			when "11000011001" => error_vector <= "0100000100000100";
			when "11000011111" => error_vector <= "0100000100000010";
			when "11000011100" => error_vector <= "0100000100000001";
			when "11111011101" => error_vector <= "0100000011000000";
			when "11110111101" => error_vector <= "0100000010100000";
			when "11110001101" => error_vector <= "0100000010010000";
			when "11110010101" => error_vector <= "0100000010001000";
			when "11110011001" => error_vector <= "0100000010000100";
			when "11110011111" => error_vector <= "0100000010000010";
			when "11110011100" => error_vector <= "0100000010000001";
			when "11101111101" => error_vector <= "0100000001100000";
			when "11101001101" => error_vector <= "0100000001010000";
			when "11101010101" => error_vector <= "0100000001001000";
			when "11101011001" => error_vector <= "0100000001000100";
			when "11101011111" => error_vector <= "0100000001000010";
			when "11101011100" => error_vector <= "0100000001000001";
			when "11100101101" => error_vector <= "0100000000110000";
			when "11100110101" => error_vector <= "0100000000101000";
			when "11100111001" => error_vector <= "0100000000100100";
			when "11100111111" => error_vector <= "0100000000100010";
			when "11100111100" => error_vector <= "0100000000100001";
			when "11100000101" => error_vector <= "0100000000011000";
			when "11100001001" => error_vector <= "0100000000010100";
			when "11100001111" => error_vector <= "0100000000010010";
			when "11100001100" => error_vector <= "0100000000010001";
			when "11100010001" => error_vector <= "0100000000001100";
			when "11100010111" => error_vector <= "0100000000001010";
			when "11100010100" => error_vector <= "0100000000001001";
			when "11100011011" => error_vector <= "0100000000000110";
			when "11100011000" => error_vector <= "0100000000000101";
			when "11100011110" => error_vector <= "0100000000000011";
			when "11100000011" => error_vector <= "0011100000000000";
			when "01001101100" => error_vector <= "0011010000000000";
			when "10001101100" => error_vector <= "0011001000000000";
			when "11101101100" => error_vector <= "0011000100000000";
			when "11011101100" => error_vector <= "0011000010000000";
			when "11000101100" => error_vector <= "0011000001000000";
			when "11001001100" => error_vector <= "0011000000100000";
			when "11001111100" => error_vector <= "0011000000010000";
			when "11001100100" => error_vector <= "0011000000001000";
			when "11001101000" => error_vector <= "0011000000000100";
			when "11001101110" => error_vector <= "0011000000000010";
			when "11001101101" => error_vector <= "0011000000000001";
			when "00110110100" => error_vector <= "0010110000000000";
			when "11110110100" => error_vector <= "0010101000000000";
			when "10010110100" => error_vector <= "0010100100000000";
			when "10100110100" => error_vector <= "0010100010000000";
			when "10111110100" => error_vector <= "0010100001000000";
			when "10110010100" => error_vector <= "0010100000100000";
			when "10110100100" => error_vector <= "0010100000010000";
			when "10110111100" => error_vector <= "0010100000001000";
			when "10110110000" => error_vector <= "0010100000000100";
			when "10110110110" => error_vector <= "0010100000000010";
			when "10110110101" => error_vector <= "0010100000000001";
			when "01011011011" => error_vector <= "0010011000000000";
			when "00111011011" => error_vector <= "0010010100000000";
			when "00001011011" => error_vector <= "0010010010000000";
			when "00010011011" => error_vector <= "0010010001000000";
			when "00011111011" => error_vector <= "0010010000100000";
			when "00011001011" => error_vector <= "0010010000010000";
			when "00011010011" => error_vector <= "0010010000001000";
			when "00011011111" => error_vector <= "0010010000000100";
			when "00011011001" => error_vector <= "0010010000000010";
			when "00011011010" => error_vector <= "0010010000000001";
			when "11111011011" => error_vector <= "0010001100000000";
			when "11001011011" => error_vector <= "0010001010000000";
			when "11010011011" => error_vector <= "0010001001000000";
			when "11011111011" => error_vector <= "0010001000100000";
			when "11011001011" => error_vector <= "0010001000010000";
			when "11011010011" => error_vector <= "0010001000001000";
			when "11011011111" => error_vector <= "0010001000000100";
			when "11011011001" => error_vector <= "0010001000000010";
			when "11011011010" => error_vector <= "0010001000000001";
			when "10101011011" => error_vector <= "0010000110000000";
			when "10110011011" => error_vector <= "0010000101000000";
			when "10111111011" => error_vector <= "0010000100100000";
			when "10111001011" => error_vector <= "0010000100010000";
			when "10111010011" => error_vector <= "0010000100001000";
			when "10111011111" => error_vector <= "0010000100000100";
			when "10111011001" => error_vector <= "0010000100000010";
			when "10111011010" => error_vector <= "0010000100000001";
			when "10000011011" => error_vector <= "0010000011000000";
			when "10001111011" => error_vector <= "0010000010100000";
			when "10001001011" => error_vector <= "0010000010010000";
			when "10001010011" => error_vector <= "0010000010001000";
			when "10001011111" => error_vector <= "0010000010000100";
			when "10001011001" => error_vector <= "0010000010000010";
			when "10001011010" => error_vector <= "0010000010000001";
			when "10010111011" => error_vector <= "0010000001100000";
			when "10010001011" => error_vector <= "0010000001010000";
			when "10010010011" => error_vector <= "0010000001001000";
			when "10010011111" => error_vector <= "0010000001000100";
			when "10010011001" => error_vector <= "0010000001000010";
			when "10010011010" => error_vector <= "0010000001000001";
			when "10011101011" => error_vector <= "0010000000110000";
			when "10011110011" => error_vector <= "0010000000101000";
			when "10011111111" => error_vector <= "0010000000100100";
			when "10011111001" => error_vector <= "0010000000100010";
			when "10011111010" => error_vector <= "0010000000100001";
			when "10011000011" => error_vector <= "0010000000011000";
			when "10011001111" => error_vector <= "0010000000010100";
			when "10011001001" => error_vector <= "0010000000010010";
			when "10011001010" => error_vector <= "0010000000010001";
			when "10011010111" => error_vector <= "0010000000001100";
			when "10011010001" => error_vector <= "0010000000001010";
			when "10011010010" => error_vector <= "0010000000001001";
			when "10011011101" => error_vector <= "0010000000000110";
			when "10011011110" => error_vector <= "0010000000000101";
			when "10011011000" => error_vector <= "0010000000000011";
			when "11111011000" => error_vector <= "0001110000000000";
			when "00111011000" => error_vector <= "0001101000000000";
			when "01011011000" => error_vector <= "0001100100000000";
			when "01101011000" => error_vector <= "0001100010000000";
			when "01110011000" => error_vector <= "0001100001000000";
			when "01111111000" => error_vector <= "0001100000100000";
			when "01111001000" => error_vector <= "0001100000010000";
			when "01111010000" => error_vector <= "0001100000001000";
			when "01111011100" => error_vector <= "0001100000000100";
			when "01111011010" => error_vector <= "0001100000000010";
			when "01111011001" => error_vector <= "0001100000000001";
			when "10010110111" => error_vector <= "0001011000000000";
			when "11110110111" => error_vector <= "0001010100000000";
			when "11000110111" => error_vector <= "0001010010000000";
			when "11011110111" => error_vector <= "0001010001000000";
			when "11010010111" => error_vector <= "0001010000100000";
			when "11010100111" => error_vector <= "0001010000010000";
			when "11010111111" => error_vector <= "0001010000001000";
			when "11010110011" => error_vector <= "0001010000000100";
			when "11010110101" => error_vector <= "0001010000000010";
			when "11010110110" => error_vector <= "0001010000000001";
			when "00110110111" => error_vector <= "0001001100000000";
			when "00000110111" => error_vector <= "0001001010000000";
			when "00011110111" => error_vector <= "0001001001000000";
			when "00010010111" => error_vector <= "0001001000100000";
			when "00010100111" => error_vector <= "0001001000010000";
			when "00010111111" => error_vector <= "0001001000001000";
			when "00010110011" => error_vector <= "0001001000000100";
			when "00010110101" => error_vector <= "0001001000000010";
			when "00010110110" => error_vector <= "0001001000000001";
			when "01100110111" => error_vector <= "0001000110000000";
			when "01111110111" => error_vector <= "0001000101000000";
			when "01110010111" => error_vector <= "0001000100100000";
			when "01110100111" => error_vector <= "0001000100010000";
			when "01110111111" => error_vector <= "0001000100001000";
			when "01110110011" => error_vector <= "0001000100000100";
			when "01110110101" => error_vector <= "0001000100000010";
			when "01110110110" => error_vector <= "0001000100000001";
			when "01001110111" => error_vector <= "0001000011000000";
			when "01000010111" => error_vector <= "0001000010100000";
			when "01000100111" => error_vector <= "0001000010010000";
			when "01000111111" => error_vector <= "0001000010001000";
			when "01000110011" => error_vector <= "0001000010000100";
			when "01000110101" => error_vector <= "0001000010000010";
			when "01000110110" => error_vector <= "0001000010000001";
			when "01011010111" => error_vector <= "0001000001100000";
			when "01011100111" => error_vector <= "0001000001010000";
			when "01011111111" => error_vector <= "0001000001001000";
			when "01011110011" => error_vector <= "0001000001000100";
			when "01011110101" => error_vector <= "0001000001000010";
			when "01011110110" => error_vector <= "0001000001000001";
			when "01010000111" => error_vector <= "0001000000110000";
			when "01010011111" => error_vector <= "0001000000101000";
			when "01010010011" => error_vector <= "0001000000100100";
			when "01010010101" => error_vector <= "0001000000100010";
			when "01010010110" => error_vector <= "0001000000100001";
			when "01010101111" => error_vector <= "0001000000011000";
			when "01010100011" => error_vector <= "0001000000010100";
			when "01010100101" => error_vector <= "0001000000010010";
			when "01010100110" => error_vector <= "0001000000010001";
			when "01010111011" => error_vector <= "0001000000001100";
			when "01010111101" => error_vector <= "0001000000001010";
			when "01010111110" => error_vector <= "0001000000001001";
			when "01010110001" => error_vector <= "0001000000000110";
			when "01010110010" => error_vector <= "0001000000000101";
			when "01010110100" => error_vector <= "0001000000000011";
			when "11101101111" => error_vector <= "0000111000000000";
			when "10001101111" => error_vector <= "0000110100000000";
			when "10111101111" => error_vector <= "0000110010000000";
			when "10100101111" => error_vector <= "0000110001000000";
			when "10101001111" => error_vector <= "0000110000100000";
			when "10101111111" => error_vector <= "0000110000010000";
			when "10101100111" => error_vector <= "0000110000001000";
			when "10101101011" => error_vector <= "0000110000000100";
			when "10101101101" => error_vector <= "0000110000000010";
			when "10101101110" => error_vector <= "0000110000000001";
			when "01001101111" => error_vector <= "0000101100000000";
			when "01111101111" => error_vector <= "0000101010000000";
			when "01100101111" => error_vector <= "0000101001000000";
			when "01101001111" => error_vector <= "0000101000100000";
			when "01101111111" => error_vector <= "0000101000010000";
			when "01101100111" => error_vector <= "0000101000001000";
			when "01101101011" => error_vector <= "0000101000000100";
			when "01101101101" => error_vector <= "0000101000000010";
			when "01101101110" => error_vector <= "0000101000000001";
			when "00011101111" => error_vector <= "0000100110000000";
			when "00000101111" => error_vector <= "0000100101000000";
			when "00001001111" => error_vector <= "0000100100100000";
			when "00001111111" => error_vector <= "0000100100010000";
			when "00001100111" => error_vector <= "0000100100001000";
			when "00001101011" => error_vector <= "0000100100000100";
			when "00001101101" => error_vector <= "0000100100000010";
			when "00001101110" => error_vector <= "0000100100000001";
			when "00110101111" => error_vector <= "0000100011000000";
			when "00111001111" => error_vector <= "0000100010100000";
			when "00111111111" => error_vector <= "0000100010010000";
			when "00111100111" => error_vector <= "0000100010001000";
			when "00111101011" => error_vector <= "0000100010000100";
			when "00111101101" => error_vector <= "0000100010000010";
			when "00111101110" => error_vector <= "0000100010000001";
			when "00100001111" => error_vector <= "0000100001100000";
			when "00100111111" => error_vector <= "0000100001010000";
			when "00100100111" => error_vector <= "0000100001001000";
			when "00100101011" => error_vector <= "0000100001000100";
			when "00100101101" => error_vector <= "0000100001000010";
			when "00100101110" => error_vector <= "0000100001000001";
			when "00101011111" => error_vector <= "0000100000110000";
			when "00101000111" => error_vector <= "0000100000101000";
			when "00101001011" => error_vector <= "0000100000100100";
			when "00101001101" => error_vector <= "0000100000100010";
			when "00101001110" => error_vector <= "0000100000100001";
			when "00101110111" => error_vector <= "0000100000011000";
			when "00101111011" => error_vector <= "0000100000010100";
			when "00101111101" => error_vector <= "0000100000010010";
			when "00101111110" => error_vector <= "0000100000010001";
			when "00101100011" => error_vector <= "0000100000001100";
			when "00101100101" => error_vector <= "0000100000001010";
			when "00101100110" => error_vector <= "0000100000001001";
			when "00101101001" => error_vector <= "0000100000000110";
			when "00101101010" => error_vector <= "0000100000000101";
			when "00101101100" => error_vector <= "0000100000000011";
			when "11100000000" => error_vector <= "0000011100000000";
			when "11010000000" => error_vector <= "0000011010000000";
			when "11001000000" => error_vector <= "0000011001000000";
			when "11000100000" => error_vector <= "0000011000100000";
			when "11000010000" => error_vector <= "0000011000010000";
			when "11000001000" => error_vector <= "0000011000001000";
			when "11000000100" => error_vector <= "0000011000000100";
			when "11000000010" => error_vector <= "0000011000000010";
			when "11000000001" => error_vector <= "0000011000000001";
			when "10110000000" => error_vector <= "0000010110000000";
			when "10101000000" => error_vector <= "0000010101000000";
			when "10100100000" => error_vector <= "0000010100100000";
			when "10100010000" => error_vector <= "0000010100010000";
			when "10100001000" => error_vector <= "0000010100001000";
			when "10100000100" => error_vector <= "0000010100000100";
			when "10100000010" => error_vector <= "0000010100000010";
			when "10100000001" => error_vector <= "0000010100000001";
			when "10011000000" => error_vector <= "0000010011000000";
			when "10010100000" => error_vector <= "0000010010100000";
			when "10010010000" => error_vector <= "0000010010010000";
			when "10010001000" => error_vector <= "0000010010001000";
			when "10010000100" => error_vector <= "0000010010000100";
			when "10010000010" => error_vector <= "0000010010000010";
			when "10010000001" => error_vector <= "0000010010000001";
			when "10001100000" => error_vector <= "0000010001100000";
			when "10001010000" => error_vector <= "0000010001010000";
			when "10001001000" => error_vector <= "0000010001001000";
			when "10001000100" => error_vector <= "0000010001000100";
			when "10001000010" => error_vector <= "0000010001000010";
			when "10001000001" => error_vector <= "0000010001000001";
			when "10000110000" => error_vector <= "0000010000110000";
			when "10000101000" => error_vector <= "0000010000101000";
			when "10000100100" => error_vector <= "0000010000100100";
			when "10000100010" => error_vector <= "0000010000100010";
			when "10000100001" => error_vector <= "0000010000100001";
			when "10000011000" => error_vector <= "0000010000011000";
			when "10000010100" => error_vector <= "0000010000010100";
			when "10000010010" => error_vector <= "0000010000010010";
			when "10000010001" => error_vector <= "0000010000010001";
			when "10000001100" => error_vector <= "0000010000001100";
			when "10000001010" => error_vector <= "0000010000001010";
			when "10000001001" => error_vector <= "0000010000001001";
			when "10000000110" => error_vector <= "0000010000000110";
			when "10000000101" => error_vector <= "0000010000000101";
			when "10000000011" => error_vector <= "0000010000000011";
			when "01110000000" => error_vector <= "0000001110000000";
			when "01101000000" => error_vector <= "0000001101000000";
			when "01100100000" => error_vector <= "0000001100100000";
			when "01100010000" => error_vector <= "0000001100010000";
			when "01100001000" => error_vector <= "0000001100001000";
			when "01100000100" => error_vector <= "0000001100000100";
			when "01100000010" => error_vector <= "0000001100000010";
			when "01100000001" => error_vector <= "0000001100000001";
			when "01011000000" => error_vector <= "0000001011000000";
			when "01010100000" => error_vector <= "0000001010100000";
			when "01010010000" => error_vector <= "0000001010010000";
			when "01010001000" => error_vector <= "0000001010001000";
			when "01010000100" => error_vector <= "0000001010000100";
			when "01010000010" => error_vector <= "0000001010000010";
			when "01010000001" => error_vector <= "0000001010000001";
			when "01001100000" => error_vector <= "0000001001100000";
			when "01001010000" => error_vector <= "0000001001010000";
			when "01001001000" => error_vector <= "0000001001001000";
			when "01001000100" => error_vector <= "0000001001000100";
			when "01001000010" => error_vector <= "0000001001000010";
			when "01001000001" => error_vector <= "0000001001000001";
			when "01000110000" => error_vector <= "0000001000110000";
			when "01000101000" => error_vector <= "0000001000101000";
			when "01000100100" => error_vector <= "0000001000100100";
			when "01000100010" => error_vector <= "0000001000100010";
			when "01000100001" => error_vector <= "0000001000100001";
			when "01000011000" => error_vector <= "0000001000011000";
			when "01000010100" => error_vector <= "0000001000010100";
			when "01000010010" => error_vector <= "0000001000010010";
			when "01000010001" => error_vector <= "0000001000010001";
			when "01000001100" => error_vector <= "0000001000001100";
			when "01000001010" => error_vector <= "0000001000001010";
			when "01000001001" => error_vector <= "0000001000001001";
			when "01000000110" => error_vector <= "0000001000000110";
			when "01000000101" => error_vector <= "0000001000000101";
			when "01000000011" => error_vector <= "0000001000000011";
			when "00111000000" => error_vector <= "0000000111000000";
			when "00110100000" => error_vector <= "0000000110100000";
			when "00110010000" => error_vector <= "0000000110010000";
			when "00110001000" => error_vector <= "0000000110001000";
			when "00110000100" => error_vector <= "0000000110000100";
			when "00110000010" => error_vector <= "0000000110000010";
			when "00110000001" => error_vector <= "0000000110000001";
			when "00101100000" => error_vector <= "0000000101100000";
			when "00101010000" => error_vector <= "0000000101010000";
			when "00101001000" => error_vector <= "0000000101001000";
			when "00101000100" => error_vector <= "0000000101000100";
			when "00101000010" => error_vector <= "0000000101000010";
			when "00101000001" => error_vector <= "0000000101000001";
			when "00100110000" => error_vector <= "0000000100110000";
			when "00100101000" => error_vector <= "0000000100101000";
			when "00100100100" => error_vector <= "0000000100100100";
			when "00100100010" => error_vector <= "0000000100100010";
			when "00100100001" => error_vector <= "0000000100100001";
			when "00100011000" => error_vector <= "0000000100011000";
			when "00100010100" => error_vector <= "0000000100010100";
			when "00100010010" => error_vector <= "0000000100010010";
			when "00100010001" => error_vector <= "0000000100010001";
			when "00100001100" => error_vector <= "0000000100001100";
			when "00100001010" => error_vector <= "0000000100001010";
			when "00100001001" => error_vector <= "0000000100001001";
			when "00100000110" => error_vector <= "0000000100000110";
			when "00100000101" => error_vector <= "0000000100000101";
			when "00100000011" => error_vector <= "0000000100000011";
			when "00011100000" => error_vector <= "0000000011100000";
			when "00011010000" => error_vector <= "0000000011010000";
			when "00011001000" => error_vector <= "0000000011001000";
			when "00011000100" => error_vector <= "0000000011000100";
			when "00011000010" => error_vector <= "0000000011000010";
			when "00011000001" => error_vector <= "0000000011000001";
			when "00010110000" => error_vector <= "0000000010110000";
			when "00010101000" => error_vector <= "0000000010101000";
			when "00010100100" => error_vector <= "0000000010100100";
			when "00010100010" => error_vector <= "0000000010100010";
			when "00010100001" => error_vector <= "0000000010100001";
			when "00010011000" => error_vector <= "0000000010011000";
			when "00010010100" => error_vector <= "0000000010010100";
			when "00010010010" => error_vector <= "0000000010010010";
			when "00010010001" => error_vector <= "0000000010010001";
			when "00010001100" => error_vector <= "0000000010001100";
			when "00010001010" => error_vector <= "0000000010001010";
			when "00010001001" => error_vector <= "0000000010001001";
			when "00010000110" => error_vector <= "0000000010000110";
			when "00010000101" => error_vector <= "0000000010000101";
			when "00010000011" => error_vector <= "0000000010000011";
			when "00001110000" => error_vector <= "0000000001110000";
			when "00001101000" => error_vector <= "0000000001101000";
			when "00001100100" => error_vector <= "0000000001100100";
			when "00001100010" => error_vector <= "0000000001100010";
			when "00001100001" => error_vector <= "0000000001100001";
			when "00001011000" => error_vector <= "0000000001011000";
			when "00001010100" => error_vector <= "0000000001010100";
			when "00001010010" => error_vector <= "0000000001010010";
			when "00001010001" => error_vector <= "0000000001010001";
			when "00001001100" => error_vector <= "0000000001001100";
			when "00001001010" => error_vector <= "0000000001001010";
			when "00001001001" => error_vector <= "0000000001001001";
			when "00001000110" => error_vector <= "0000000001000110";
			when "00001000101" => error_vector <= "0000000001000101";
			when "00001000011" => error_vector <= "0000000001000011";
			when "00000111000" => error_vector <= "0000000000111000";
			when "00000110100" => error_vector <= "0000000000110100";
			when "00000110010" => error_vector <= "0000000000110010";
			when "00000110001" => error_vector <= "0000000000110001";
			when "00000101100" => error_vector <= "0000000000101100";
			when "00000101010" => error_vector <= "0000000000101010";
			when "00000101001" => error_vector <= "0000000000101001";
			when "00000100110" => error_vector <= "0000000000100110";
			when "00000100101" => error_vector <= "0000000000100101";
			when "00000100011" => error_vector <= "0000000000100011";
			when "00000011100" => error_vector <= "0000000000011100";
			when "00000011010" => error_vector <= "0000000000011010";
			when "00000011001" => error_vector <= "0000000000011001";
			when "00000010110" => error_vector <= "0000000000010110";
			when "00000010101" => error_vector <= "0000000000010101";
			when "00000010011" => error_vector <= "0000000000010011";
			when "00000001110" => error_vector <= "0000000000001110";
			when "00000001101" => error_vector <= "0000000000001101";
			when "00000001011" => error_vector <= "0000000000001011";
			when "00000000111" => error_vector <= "0000000000000111";
			when others	=> error_vector <= "0000000000000000";
		end case check_syndromes;
	end process;
end corr; -- syndrome_correction.