module reg1000 ( in, clk, rst, out );
	input[31:0] in;
	input clk;
	input rst;
	output[31:0] out;

	wire [31:0] r0_out;
	wire [31:0] r1_out;
	wire [31:0] r2_out;
	wire [31:0] r3_out;
	wire [31:0] r4_out;
	wire [31:0] r5_out;
	wire [31:0] r6_out;
	wire [31:0] r7_out;
	wire [31:0] r8_out;
	wire [31:0] r9_out;
	wire [31:0] r10_out;
	wire [31:0] r11_out;
	wire [31:0] r12_out;
	wire [31:0] r13_out;
	wire [31:0] r14_out;
	wire [31:0] r15_out;
	wire [31:0] r16_out;
	wire [31:0] r17_out;
	wire [31:0] r18_out;
	wire [31:0] r19_out;
	wire [31:0] r20_out;
	wire [31:0] r21_out;
	wire [31:0] r22_out;
	wire [31:0] r23_out;
	wire [31:0] r24_out;
	wire [31:0] r25_out;
	wire [31:0] r26_out;
	wire [31:0] r27_out;
	wire [31:0] r28_out;
	wire [31:0] r29_out;
	wire [31:0] r30_out;
	wire [31:0] r31_out;
	wire [31:0] r32_out;
	wire [31:0] r33_out;
	wire [31:0] r34_out;
	wire [31:0] r35_out;
	wire [31:0] r36_out;
	wire [31:0] r37_out;
	wire [31:0] r38_out;
	wire [31:0] r39_out;
	wire [31:0] r40_out;
	wire [31:0] r41_out;
	wire [31:0] r42_out;
	wire [31:0] r43_out;
	wire [31:0] r44_out;
	wire [31:0] r45_out;
	wire [31:0] r46_out;
	wire [31:0] r47_out;
	wire [31:0] r48_out;
	wire [31:0] r49_out;
	wire [31:0] r50_out;
	wire [31:0] r51_out;
	wire [31:0] r52_out;
	wire [31:0] r53_out;
	wire [31:0] r54_out;
	wire [31:0] r55_out;
	wire [31:0] r56_out;
	wire [31:0] r57_out;
	wire [31:0] r58_out;
	wire [31:0] r59_out;
	wire [31:0] r60_out;
	wire [31:0] r61_out;
	wire [31:0] r62_out;
	wire [31:0] r63_out;
	wire [31:0] r64_out;
	wire [31:0] r65_out;
	wire [31:0] r66_out;
	wire [31:0] r67_out;
	wire [31:0] r68_out;
	wire [31:0] r69_out;
	wire [31:0] r70_out;
	wire [31:0] r71_out;
	wire [31:0] r72_out;
	wire [31:0] r73_out;
	wire [31:0] r74_out;
	wire [31:0] r75_out;
	wire [31:0] r76_out;
	wire [31:0] r77_out;
	wire [31:0] r78_out;
	wire [31:0] r79_out;
	wire [31:0] r80_out;
	wire [31:0] r81_out;
	wire [31:0] r82_out;
	wire [31:0] r83_out;
	wire [31:0] r84_out;
	wire [31:0] r85_out;
	wire [31:0] r86_out;
	wire [31:0] r87_out;
	wire [31:0] r88_out;
	wire [31:0] r89_out;
	wire [31:0] r90_out;
	wire [31:0] r91_out;
	wire [31:0] r92_out;
	wire [31:0] r93_out;
	wire [31:0] r94_out;
	wire [31:0] r95_out;
	wire [31:0] r96_out;
	wire [31:0] r97_out;
	wire [31:0] r98_out;
	wire [31:0] r99_out;
	wire [31:0] r100_out;
	wire [31:0] r101_out;
	wire [31:0] r102_out;
	wire [31:0] r103_out;
	wire [31:0] r104_out;
	wire [31:0] r105_out;
	wire [31:0] r106_out;
	wire [31:0] r107_out;
	wire [31:0] r108_out;
	wire [31:0] r109_out;
	wire [31:0] r110_out;
	wire [31:0] r111_out;
	wire [31:0] r112_out;
	wire [31:0] r113_out;
	wire [31:0] r114_out;
	wire [31:0] r115_out;
	wire [31:0] r116_out;
	wire [31:0] r117_out;
	wire [31:0] r118_out;
	wire [31:0] r119_out;
	wire [31:0] r120_out;
	wire [31:0] r121_out;
	wire [31:0] r122_out;
	wire [31:0] r123_out;
	wire [31:0] r124_out;
	wire [31:0] r125_out;
	wire [31:0] r126_out;
	wire [31:0] r127_out;
	wire [31:0] r128_out;
	wire [31:0] r129_out;
	wire [31:0] r130_out;
	wire [31:0] r131_out;
	wire [31:0] r132_out;
	wire [31:0] r133_out;
	wire [31:0] r134_out;
	wire [31:0] r135_out;
	wire [31:0] r136_out;
	wire [31:0] r137_out;
	wire [31:0] r138_out;
	wire [31:0] r139_out;
	wire [31:0] r140_out;
	wire [31:0] r141_out;
	wire [31:0] r142_out;
	wire [31:0] r143_out;
	wire [31:0] r144_out;
	wire [31:0] r145_out;
	wire [31:0] r146_out;
	wire [31:0] r147_out;
	wire [31:0] r148_out;
	wire [31:0] r149_out;
	wire [31:0] r150_out;
	wire [31:0] r151_out;
	wire [31:0] r152_out;
	wire [31:0] r153_out;
	wire [31:0] r154_out;
	wire [31:0] r155_out;
	wire [31:0] r156_out;
	wire [31:0] r157_out;
	wire [31:0] r158_out;
	wire [31:0] r159_out;
	wire [31:0] r160_out;
	wire [31:0] r161_out;
	wire [31:0] r162_out;
	wire [31:0] r163_out;
	wire [31:0] r164_out;
	wire [31:0] r165_out;
	wire [31:0] r166_out;
	wire [31:0] r167_out;
	wire [31:0] r168_out;
	wire [31:0] r169_out;
	wire [31:0] r170_out;
	wire [31:0] r171_out;
	wire [31:0] r172_out;
	wire [31:0] r173_out;
	wire [31:0] r174_out;
	wire [31:0] r175_out;
	wire [31:0] r176_out;
	wire [31:0] r177_out;
	wire [31:0] r178_out;
	wire [31:0] r179_out;
	wire [31:0] r180_out;
	wire [31:0] r181_out;
	wire [31:0] r182_out;
	wire [31:0] r183_out;
	wire [31:0] r184_out;
	wire [31:0] r185_out;
	wire [31:0] r186_out;
	wire [31:0] r187_out;
	wire [31:0] r188_out;
	wire [31:0] r189_out;
	wire [31:0] r190_out;
	wire [31:0] r191_out;
	wire [31:0] r192_out;
	wire [31:0] r193_out;
	wire [31:0] r194_out;
	wire [31:0] r195_out;
	wire [31:0] r196_out;
	wire [31:0] r197_out;
	wire [31:0] r198_out;
	wire [31:0] r199_out;
	wire [31:0] r200_out;
	wire [31:0] r201_out;
	wire [31:0] r202_out;
	wire [31:0] r203_out;
	wire [31:0] r204_out;
	wire [31:0] r205_out;
	wire [31:0] r206_out;
	wire [31:0] r207_out;
	wire [31:0] r208_out;
	wire [31:0] r209_out;
	wire [31:0] r210_out;
	wire [31:0] r211_out;
	wire [31:0] r212_out;
	wire [31:0] r213_out;
	wire [31:0] r214_out;
	wire [31:0] r215_out;
	wire [31:0] r216_out;
	wire [31:0] r217_out;
	wire [31:0] r218_out;
	wire [31:0] r219_out;
	wire [31:0] r220_out;
	wire [31:0] r221_out;
	wire [31:0] r222_out;
	wire [31:0] r223_out;
	wire [31:0] r224_out;
	wire [31:0] r225_out;
	wire [31:0] r226_out;
	wire [31:0] r227_out;
	wire [31:0] r228_out;
	wire [31:0] r229_out;
	wire [31:0] r230_out;
	wire [31:0] r231_out;
	wire [31:0] r232_out;
	wire [31:0] r233_out;
	wire [31:0] r234_out;
	wire [31:0] r235_out;
	wire [31:0] r236_out;
	wire [31:0] r237_out;
	wire [31:0] r238_out;
	wire [31:0] r239_out;
	wire [31:0] r240_out;
	wire [31:0] r241_out;
	wire [31:0] r242_out;
	wire [31:0] r243_out;
	wire [31:0] r244_out;
	wire [31:0] r245_out;
	wire [31:0] r246_out;
	wire [31:0] r247_out;
	wire [31:0] r248_out;
	wire [31:0] r249_out;
	wire [31:0] r250_out;
	wire [31:0] r251_out;
	wire [31:0] r252_out;
	wire [31:0] r253_out;
	wire [31:0] r254_out;
	wire [31:0] r255_out;
	wire [31:0] r256_out;
	wire [31:0] r257_out;
	wire [31:0] r258_out;
	wire [31:0] r259_out;
	wire [31:0] r260_out;
	wire [31:0] r261_out;
	wire [31:0] r262_out;
	wire [31:0] r263_out;
	wire [31:0] r264_out;
	wire [31:0] r265_out;
	wire [31:0] r266_out;
	wire [31:0] r267_out;
	wire [31:0] r268_out;
	wire [31:0] r269_out;
	wire [31:0] r270_out;
	wire [31:0] r271_out;
	wire [31:0] r272_out;
	wire [31:0] r273_out;
	wire [31:0] r274_out;
	wire [31:0] r275_out;
	wire [31:0] r276_out;
	wire [31:0] r277_out;
	wire [31:0] r278_out;
	wire [31:0] r279_out;
	wire [31:0] r280_out;
	wire [31:0] r281_out;
	wire [31:0] r282_out;
	wire [31:0] r283_out;
	wire [31:0] r284_out;
	wire [31:0] r285_out;
	wire [31:0] r286_out;
	wire [31:0] r287_out;
	wire [31:0] r288_out;
	wire [31:0] r289_out;
	wire [31:0] r290_out;
	wire [31:0] r291_out;
	wire [31:0] r292_out;
	wire [31:0] r293_out;
	wire [31:0] r294_out;
	wire [31:0] r295_out;
	wire [31:0] r296_out;
	wire [31:0] r297_out;
	wire [31:0] r298_out;
	wire [31:0] r299_out;
	wire [31:0] r300_out;
	wire [31:0] r301_out;
	wire [31:0] r302_out;
	wire [31:0] r303_out;
	wire [31:0] r304_out;
	wire [31:0] r305_out;
	wire [31:0] r306_out;
	wire [31:0] r307_out;
	wire [31:0] r308_out;
	wire [31:0] r309_out;
	wire [31:0] r310_out;
	wire [31:0] r311_out;
	wire [31:0] r312_out;
	wire [31:0] r313_out;
	wire [31:0] r314_out;
	wire [31:0] r315_out;
	wire [31:0] r316_out;
	wire [31:0] r317_out;
	wire [31:0] r318_out;
	wire [31:0] r319_out;
	wire [31:0] r320_out;
	wire [31:0] r321_out;
	wire [31:0] r322_out;
	wire [31:0] r323_out;
	wire [31:0] r324_out;
	wire [31:0] r325_out;
	wire [31:0] r326_out;
	wire [31:0] r327_out;
	wire [31:0] r328_out;
	wire [31:0] r329_out;
	wire [31:0] r330_out;
	wire [31:0] r331_out;
	wire [31:0] r332_out;
	wire [31:0] r333_out;
	wire [31:0] r334_out;
	wire [31:0] r335_out;
	wire [31:0] r336_out;
	wire [31:0] r337_out;
	wire [31:0] r338_out;
	wire [31:0] r339_out;
	wire [31:0] r340_out;
	wire [31:0] r341_out;
	wire [31:0] r342_out;
	wire [31:0] r343_out;
	wire [31:0] r344_out;
	wire [31:0] r345_out;
	wire [31:0] r346_out;
	wire [31:0] r347_out;
	wire [31:0] r348_out;
	wire [31:0] r349_out;
	wire [31:0] r350_out;
	wire [31:0] r351_out;
	wire [31:0] r352_out;
	wire [31:0] r353_out;
	wire [31:0] r354_out;
	wire [31:0] r355_out;
	wire [31:0] r356_out;
	wire [31:0] r357_out;
	wire [31:0] r358_out;
	wire [31:0] r359_out;
	wire [31:0] r360_out;
	wire [31:0] r361_out;
	wire [31:0] r362_out;
	wire [31:0] r363_out;
	wire [31:0] r364_out;
	wire [31:0] r365_out;
	wire [31:0] r366_out;
	wire [31:0] r367_out;
	wire [31:0] r368_out;
	wire [31:0] r369_out;
	wire [31:0] r370_out;
	wire [31:0] r371_out;
	wire [31:0] r372_out;
	wire [31:0] r373_out;
	wire [31:0] r374_out;
	wire [31:0] r375_out;
	wire [31:0] r376_out;
	wire [31:0] r377_out;
	wire [31:0] r378_out;
	wire [31:0] r379_out;
	wire [31:0] r380_out;
	wire [31:0] r381_out;
	wire [31:0] r382_out;
	wire [31:0] r383_out;
	wire [31:0] r384_out;
	wire [31:0] r385_out;
	wire [31:0] r386_out;
	wire [31:0] r387_out;
	wire [31:0] r388_out;
	wire [31:0] r389_out;
	wire [31:0] r390_out;
	wire [31:0] r391_out;
	wire [31:0] r392_out;
	wire [31:0] r393_out;
	wire [31:0] r394_out;
	wire [31:0] r395_out;
	wire [31:0] r396_out;
	wire [31:0] r397_out;
	wire [31:0] r398_out;
	wire [31:0] r399_out;
	wire [31:0] r400_out;
	wire [31:0] r401_out;
	wire [31:0] r402_out;
	wire [31:0] r403_out;
	wire [31:0] r404_out;
	wire [31:0] r405_out;
	wire [31:0] r406_out;
	wire [31:0] r407_out;
	wire [31:0] r408_out;
	wire [31:0] r409_out;
	wire [31:0] r410_out;
	wire [31:0] r411_out;
	wire [31:0] r412_out;
	wire [31:0] r413_out;
	wire [31:0] r414_out;
	wire [31:0] r415_out;
	wire [31:0] r416_out;
	wire [31:0] r417_out;
	wire [31:0] r418_out;
	wire [31:0] r419_out;
	wire [31:0] r420_out;
	wire [31:0] r421_out;
	wire [31:0] r422_out;
	wire [31:0] r423_out;
	wire [31:0] r424_out;
	wire [31:0] r425_out;
	wire [31:0] r426_out;
	wire [31:0] r427_out;
	wire [31:0] r428_out;
	wire [31:0] r429_out;
	wire [31:0] r430_out;
	wire [31:0] r431_out;
	wire [31:0] r432_out;
	wire [31:0] r433_out;
	wire [31:0] r434_out;
	wire [31:0] r435_out;
	wire [31:0] r436_out;
	wire [31:0] r437_out;
	wire [31:0] r438_out;
	wire [31:0] r439_out;
	wire [31:0] r440_out;
	wire [31:0] r441_out;
	wire [31:0] r442_out;
	wire [31:0] r443_out;
	wire [31:0] r444_out;
	wire [31:0] r445_out;
	wire [31:0] r446_out;
	wire [31:0] r447_out;
	wire [31:0] r448_out;
	wire [31:0] r449_out;
	wire [31:0] r450_out;
	wire [31:0] r451_out;
	wire [31:0] r452_out;
	wire [31:0] r453_out;
	wire [31:0] r454_out;
	wire [31:0] r455_out;
	wire [31:0] r456_out;
	wire [31:0] r457_out;
	wire [31:0] r458_out;
	wire [31:0] r459_out;
	wire [31:0] r460_out;
	wire [31:0] r461_out;
	wire [31:0] r462_out;
	wire [31:0] r463_out;
	wire [31:0] r464_out;
	wire [31:0] r465_out;
	wire [31:0] r466_out;
	wire [31:0] r467_out;
	wire [31:0] r468_out;
	wire [31:0] r469_out;
	wire [31:0] r470_out;
	wire [31:0] r471_out;
	wire [31:0] r472_out;
	wire [31:0] r473_out;
	wire [31:0] r474_out;
	wire [31:0] r475_out;
	wire [31:0] r476_out;
	wire [31:0] r477_out;
	wire [31:0] r478_out;
	wire [31:0] r479_out;
	wire [31:0] r480_out;
	wire [31:0] r481_out;
	wire [31:0] r482_out;
	wire [31:0] r483_out;
	wire [31:0] r484_out;
	wire [31:0] r485_out;
	wire [31:0] r486_out;
	wire [31:0] r487_out;
	wire [31:0] r488_out;
	wire [31:0] r489_out;
	wire [31:0] r490_out;
	wire [31:0] r491_out;
	wire [31:0] r492_out;
	wire [31:0] r493_out;
	wire [31:0] r494_out;
	wire [31:0] r495_out;
	wire [31:0] r496_out;
	wire [31:0] r497_out;
	wire [31:0] r498_out;
	wire [31:0] r499_out;
	wire [31:0] r500_out;
	wire [31:0] r501_out;
	wire [31:0] r502_out;
	wire [31:0] r503_out;
	wire [31:0] r504_out;
	wire [31:0] r505_out;
	wire [31:0] r506_out;
	wire [31:0] r507_out;
	wire [31:0] r508_out;
	wire [31:0] r509_out;
	wire [31:0] r510_out;
	wire [31:0] r511_out;
	wire [31:0] r512_out;
	wire [31:0] r513_out;
	wire [31:0] r514_out;
	wire [31:0] r515_out;
	wire [31:0] r516_out;
	wire [31:0] r517_out;
	wire [31:0] r518_out;
	wire [31:0] r519_out;
	wire [31:0] r520_out;
	wire [31:0] r521_out;
	wire [31:0] r522_out;
	wire [31:0] r523_out;
	wire [31:0] r524_out;
	wire [31:0] r525_out;
	wire [31:0] r526_out;
	wire [31:0] r527_out;
	wire [31:0] r528_out;
	wire [31:0] r529_out;
	wire [31:0] r530_out;
	wire [31:0] r531_out;
	wire [31:0] r532_out;
	wire [31:0] r533_out;
	wire [31:0] r534_out;
	wire [31:0] r535_out;
	wire [31:0] r536_out;
	wire [31:0] r537_out;
	wire [31:0] r538_out;
	wire [31:0] r539_out;
	wire [31:0] r540_out;
	wire [31:0] r541_out;
	wire [31:0] r542_out;
	wire [31:0] r543_out;
	wire [31:0] r544_out;
	wire [31:0] r545_out;
	wire [31:0] r546_out;
	wire [31:0] r547_out;
	wire [31:0] r548_out;
	wire [31:0] r549_out;
	wire [31:0] r550_out;
	wire [31:0] r551_out;
	wire [31:0] r552_out;
	wire [31:0] r553_out;
	wire [31:0] r554_out;
	wire [31:0] r555_out;
	wire [31:0] r556_out;
	wire [31:0] r557_out;
	wire [31:0] r558_out;
	wire [31:0] r559_out;
	wire [31:0] r560_out;
	wire [31:0] r561_out;
	wire [31:0] r562_out;
	wire [31:0] r563_out;
	wire [31:0] r564_out;
	wire [31:0] r565_out;
	wire [31:0] r566_out;
	wire [31:0] r567_out;
	wire [31:0] r568_out;
	wire [31:0] r569_out;
	wire [31:0] r570_out;
	wire [31:0] r571_out;
	wire [31:0] r572_out;
	wire [31:0] r573_out;
	wire [31:0] r574_out;
	wire [31:0] r575_out;
	wire [31:0] r576_out;
	wire [31:0] r577_out;
	wire [31:0] r578_out;
	wire [31:0] r579_out;
	wire [31:0] r580_out;
	wire [31:0] r581_out;
	wire [31:0] r582_out;
	wire [31:0] r583_out;
	wire [31:0] r584_out;
	wire [31:0] r585_out;
	wire [31:0] r586_out;
	wire [31:0] r587_out;
	wire [31:0] r588_out;
	wire [31:0] r589_out;
	wire [31:0] r590_out;
	wire [31:0] r591_out;
	wire [31:0] r592_out;
	wire [31:0] r593_out;
	wire [31:0] r594_out;
	wire [31:0] r595_out;
	wire [31:0] r596_out;
	wire [31:0] r597_out;
	wire [31:0] r598_out;
	wire [31:0] r599_out;
	wire [31:0] r600_out;
	wire [31:0] r601_out;
	wire [31:0] r602_out;
	wire [31:0] r603_out;
	wire [31:0] r604_out;
	wire [31:0] r605_out;
	wire [31:0] r606_out;
	wire [31:0] r607_out;
	wire [31:0] r608_out;
	wire [31:0] r609_out;
	wire [31:0] r610_out;
	wire [31:0] r611_out;
	wire [31:0] r612_out;
	wire [31:0] r613_out;
	wire [31:0] r614_out;
	wire [31:0] r615_out;
	wire [31:0] r616_out;
	wire [31:0] r617_out;
	wire [31:0] r618_out;
	wire [31:0] r619_out;
	wire [31:0] r620_out;
	wire [31:0] r621_out;
	wire [31:0] r622_out;
	wire [31:0] r623_out;
	wire [31:0] r624_out;
	wire [31:0] r625_out;
	wire [31:0] r626_out;
	wire [31:0] r627_out;
	wire [31:0] r628_out;
	wire [31:0] r629_out;
	wire [31:0] r630_out;
	wire [31:0] r631_out;
	wire [31:0] r632_out;
	wire [31:0] r633_out;
	wire [31:0] r634_out;
	wire [31:0] r635_out;
	wire [31:0] r636_out;
	wire [31:0] r637_out;
	wire [31:0] r638_out;
	wire [31:0] r639_out;
	wire [31:0] r640_out;
	wire [31:0] r641_out;
	wire [31:0] r642_out;
	wire [31:0] r643_out;
	wire [31:0] r644_out;
	wire [31:0] r645_out;
	wire [31:0] r646_out;
	wire [31:0] r647_out;
	wire [31:0] r648_out;
	wire [31:0] r649_out;
	wire [31:0] r650_out;
	wire [31:0] r651_out;
	wire [31:0] r652_out;
	wire [31:0] r653_out;
	wire [31:0] r654_out;
	wire [31:0] r655_out;
	wire [31:0] r656_out;
	wire [31:0] r657_out;
	wire [31:0] r658_out;
	wire [31:0] r659_out;
	wire [31:0] r660_out;
	wire [31:0] r661_out;
	wire [31:0] r662_out;
	wire [31:0] r663_out;
	wire [31:0] r664_out;
	wire [31:0] r665_out;
	wire [31:0] r666_out;
	wire [31:0] r667_out;
	wire [31:0] r668_out;
	wire [31:0] r669_out;
	wire [31:0] r670_out;
	wire [31:0] r671_out;
	wire [31:0] r672_out;
	wire [31:0] r673_out;
	wire [31:0] r674_out;
	wire [31:0] r675_out;
	wire [31:0] r676_out;
	wire [31:0] r677_out;
	wire [31:0] r678_out;
	wire [31:0] r679_out;
	wire [31:0] r680_out;
	wire [31:0] r681_out;
	wire [31:0] r682_out;
	wire [31:0] r683_out;
	wire [31:0] r684_out;
	wire [31:0] r685_out;
	wire [31:0] r686_out;
	wire [31:0] r687_out;
	wire [31:0] r688_out;
	wire [31:0] r689_out;
	wire [31:0] r690_out;
	wire [31:0] r691_out;
	wire [31:0] r692_out;
	wire [31:0] r693_out;
	wire [31:0] r694_out;
	wire [31:0] r695_out;
	wire [31:0] r696_out;
	wire [31:0] r697_out;
	wire [31:0] r698_out;
	wire [31:0] r699_out;
	wire [31:0] r700_out;
	wire [31:0] r701_out;
	wire [31:0] r702_out;
	wire [31:0] r703_out;
	wire [31:0] r704_out;
	wire [31:0] r705_out;
	wire [31:0] r706_out;
	wire [31:0] r707_out;
	wire [31:0] r708_out;
	wire [31:0] r709_out;
	wire [31:0] r710_out;
	wire [31:0] r711_out;
	wire [31:0] r712_out;
	wire [31:0] r713_out;
	wire [31:0] r714_out;
	wire [31:0] r715_out;
	wire [31:0] r716_out;
	wire [31:0] r717_out;
	wire [31:0] r718_out;
	wire [31:0] r719_out;
	wire [31:0] r720_out;
	wire [31:0] r721_out;
	wire [31:0] r722_out;
	wire [31:0] r723_out;
	wire [31:0] r724_out;
	wire [31:0] r725_out;
	wire [31:0] r726_out;
	wire [31:0] r727_out;
	wire [31:0] r728_out;
	wire [31:0] r729_out;
	wire [31:0] r730_out;
	wire [31:0] r731_out;
	wire [31:0] r732_out;
	wire [31:0] r733_out;
	wire [31:0] r734_out;
	wire [31:0] r735_out;
	wire [31:0] r736_out;
	wire [31:0] r737_out;
	wire [31:0] r738_out;
	wire [31:0] r739_out;
	wire [31:0] r740_out;
	wire [31:0] r741_out;
	wire [31:0] r742_out;
	wire [31:0] r743_out;
	wire [31:0] r744_out;
	wire [31:0] r745_out;
	wire [31:0] r746_out;
	wire [31:0] r747_out;
	wire [31:0] r748_out;
	wire [31:0] r749_out;
	wire [31:0] r750_out;
	wire [31:0] r751_out;
	wire [31:0] r752_out;
	wire [31:0] r753_out;
	wire [31:0] r754_out;
	wire [31:0] r755_out;
	wire [31:0] r756_out;
	wire [31:0] r757_out;
	wire [31:0] r758_out;
	wire [31:0] r759_out;
	wire [31:0] r760_out;
	wire [31:0] r761_out;
	wire [31:0] r762_out;
	wire [31:0] r763_out;
	wire [31:0] r764_out;
	wire [31:0] r765_out;
	wire [31:0] r766_out;
	wire [31:0] r767_out;
	wire [31:0] r768_out;
	wire [31:0] r769_out;
	wire [31:0] r770_out;
	wire [31:0] r771_out;
	wire [31:0] r772_out;
	wire [31:0] r773_out;
	wire [31:0] r774_out;
	wire [31:0] r775_out;
	wire [31:0] r776_out;
	wire [31:0] r777_out;
	wire [31:0] r778_out;
	wire [31:0] r779_out;
	wire [31:0] r780_out;
	wire [31:0] r781_out;
	wire [31:0] r782_out;
	wire [31:0] r783_out;
	wire [31:0] r784_out;
	wire [31:0] r785_out;
	wire [31:0] r786_out;
	wire [31:0] r787_out;
	wire [31:0] r788_out;
	wire [31:0] r789_out;
	wire [31:0] r790_out;
	wire [31:0] r791_out;
	wire [31:0] r792_out;
	wire [31:0] r793_out;
	wire [31:0] r794_out;
	wire [31:0] r795_out;
	wire [31:0] r796_out;
	wire [31:0] r797_out;
	wire [31:0] r798_out;
	wire [31:0] r799_out;
	wire [31:0] r800_out;
	wire [31:0] r801_out;
	wire [31:0] r802_out;
	wire [31:0] r803_out;
	wire [31:0] r804_out;
	wire [31:0] r805_out;
	wire [31:0] r806_out;
	wire [31:0] r807_out;
	wire [31:0] r808_out;
	wire [31:0] r809_out;
	wire [31:0] r810_out;
	wire [31:0] r811_out;
	wire [31:0] r812_out;
	wire [31:0] r813_out;
	wire [31:0] r814_out;
	wire [31:0] r815_out;
	wire [31:0] r816_out;
	wire [31:0] r817_out;
	wire [31:0] r818_out;
	wire [31:0] r819_out;
	wire [31:0] r820_out;
	wire [31:0] r821_out;
	wire [31:0] r822_out;
	wire [31:0] r823_out;
	wire [31:0] r824_out;
	wire [31:0] r825_out;
	wire [31:0] r826_out;
	wire [31:0] r827_out;
	wire [31:0] r828_out;
	wire [31:0] r829_out;
	wire [31:0] r830_out;
	wire [31:0] r831_out;
	wire [31:0] r832_out;
	wire [31:0] r833_out;
	wire [31:0] r834_out;
	wire [31:0] r835_out;
	wire [31:0] r836_out;
	wire [31:0] r837_out;
	wire [31:0] r838_out;
	wire [31:0] r839_out;
	wire [31:0] r840_out;
	wire [31:0] r841_out;
	wire [31:0] r842_out;
	wire [31:0] r843_out;
	wire [31:0] r844_out;
	wire [31:0] r845_out;
	wire [31:0] r846_out;
	wire [31:0] r847_out;
	wire [31:0] r848_out;
	wire [31:0] r849_out;
	wire [31:0] r850_out;
	wire [31:0] r851_out;
	wire [31:0] r852_out;
	wire [31:0] r853_out;
	wire [31:0] r854_out;
	wire [31:0] r855_out;
	wire [31:0] r856_out;
	wire [31:0] r857_out;
	wire [31:0] r858_out;
	wire [31:0] r859_out;
	wire [31:0] r860_out;
	wire [31:0] r861_out;
	wire [31:0] r862_out;
	wire [31:0] r863_out;
	wire [31:0] r864_out;
	wire [31:0] r865_out;
	wire [31:0] r866_out;
	wire [31:0] r867_out;
	wire [31:0] r868_out;
	wire [31:0] r869_out;
	wire [31:0] r870_out;
	wire [31:0] r871_out;
	wire [31:0] r872_out;
	wire [31:0] r873_out;
	wire [31:0] r874_out;
	wire [31:0] r875_out;
	wire [31:0] r876_out;
	wire [31:0] r877_out;
	wire [31:0] r878_out;
	wire [31:0] r879_out;
	wire [31:0] r880_out;
	wire [31:0] r881_out;
	wire [31:0] r882_out;
	wire [31:0] r883_out;
	wire [31:0] r884_out;
	wire [31:0] r885_out;
	wire [31:0] r886_out;
	wire [31:0] r887_out;
	wire [31:0] r888_out;
	wire [31:0] r889_out;
	wire [31:0] r890_out;
	wire [31:0] r891_out;
	wire [31:0] r892_out;
	wire [31:0] r893_out;
	wire [31:0] r894_out;
	wire [31:0] r895_out;
	wire [31:0] r896_out;
	wire [31:0] r897_out;
	wire [31:0] r898_out;
	wire [31:0] r899_out;
	wire [31:0] r900_out;
	wire [31:0] r901_out;
	wire [31:0] r902_out;
	wire [31:0] r903_out;
	wire [31:0] r904_out;
	wire [31:0] r905_out;
	wire [31:0] r906_out;
	wire [31:0] r907_out;
	wire [31:0] r908_out;
	wire [31:0] r909_out;
	wire [31:0] r910_out;
	wire [31:0] r911_out;
	wire [31:0] r912_out;
	wire [31:0] r913_out;
	wire [31:0] r914_out;
	wire [31:0] r915_out;
	wire [31:0] r916_out;
	wire [31:0] r917_out;
	wire [31:0] r918_out;
	wire [31:0] r919_out;
	wire [31:0] r920_out;
	wire [31:0] r921_out;
	wire [31:0] r922_out;
	wire [31:0] r923_out;
	wire [31:0] r924_out;
	wire [31:0] r925_out;
	wire [31:0] r926_out;
	wire [31:0] r927_out;
	wire [31:0] r928_out;
	wire [31:0] r929_out;
	wire [31:0] r930_out;
	wire [31:0] r931_out;
	wire [31:0] r932_out;
	wire [31:0] r933_out;
	wire [31:0] r934_out;
	wire [31:0] r935_out;
	wire [31:0] r936_out;
	wire [31:0] r937_out;
	wire [31:0] r938_out;
	wire [31:0] r939_out;
	wire [31:0] r940_out;
	wire [31:0] r941_out;
	wire [31:0] r942_out;
	wire [31:0] r943_out;
	wire [31:0] r944_out;
	wire [31:0] r945_out;
	wire [31:0] r946_out;
	wire [31:0] r947_out;
	wire [31:0] r948_out;
	wire [31:0] r949_out;
	wire [31:0] r950_out;
	wire [31:0] r951_out;
	wire [31:0] r952_out;
	wire [31:0] r953_out;
	wire [31:0] r954_out;
	wire [31:0] r955_out;
	wire [31:0] r956_out;
	wire [31:0] r957_out;
	wire [31:0] r958_out;
	wire [31:0] r959_out;
	wire [31:0] r960_out;
	wire [31:0] r961_out;
	wire [31:0] r962_out;
	wire [31:0] r963_out;
	wire [31:0] r964_out;
	wire [31:0] r965_out;
	wire [31:0] r966_out;
	wire [31:0] r967_out;
	wire [31:0] r968_out;
	wire [31:0] r969_out;
	wire [31:0] r970_out;
	wire [31:0] r971_out;
	wire [31:0] r972_out;
	wire [31:0] r973_out;
	wire [31:0] r974_out;
	wire [31:0] r975_out;
	wire [31:0] r976_out;
	wire [31:0] r977_out;
	wire [31:0] r978_out;
	wire [31:0] r979_out;
	wire [31:0] r980_out;
	wire [31:0] r981_out;
	wire [31:0] r982_out;
	wire [31:0] r983_out;
	wire [31:0] r984_out;
	wire [31:0] r985_out;
	wire [31:0] r986_out;
	wire [31:0] r987_out;
	wire [31:0] r988_out;
	wire [31:0] r989_out;
	wire [31:0] r990_out;
	wire [31:0] r991_out;
	wire [31:0] r992_out;
	wire [31:0] r993_out;
	wire [31:0] r994_out;
	wire [31:0] r995_out;
	wire [31:0] r996_out;
	wire [31:0] r997_out;
	wire [31:0] r998_out;
	wire [31:0] r999_out;

	reg32 r0 (rst, clk, in, r0_out);
	reg32 r1 (rst, clk, r0_out, r1_out);
	reg32 r2 (rst, clk, r1_out, r2_out);
	reg32 r3 (rst, clk, r2_out, r3_out);
	reg32 r4 (rst, clk, r3_out, r4_out);
	reg32 r5 (rst, clk, r4_out, r5_out);
	reg32 r6 (rst, clk, r5_out, r6_out);
	reg32 r7 (rst, clk, r6_out, r7_out);
	reg32 r8 (rst, clk, r7_out, r8_out);
	reg32 r9 (rst, clk, r8_out, r9_out);
	reg32 r10 (rst, clk, r9_out, r10_out);
	reg32 r11 (rst, clk, r10_out, r11_out);
	reg32 r12 (rst, clk, r11_out, r12_out);
	reg32 r13 (rst, clk, r12_out, r13_out);
	reg32 r14 (rst, clk, r13_out, r14_out);
	reg32 r15 (rst, clk, r14_out, r15_out);
	reg32 r16 (rst, clk, r15_out, r16_out);
	reg32 r17 (rst, clk, r16_out, r17_out);
	reg32 r18 (rst, clk, r17_out, r18_out);
	reg32 r19 (rst, clk, r18_out, r19_out);
	reg32 r20 (rst, clk, r19_out, r20_out);
	reg32 r21 (rst, clk, r20_out, r21_out);
	reg32 r22 (rst, clk, r21_out, r22_out);
	reg32 r23 (rst, clk, r22_out, r23_out);
	reg32 r24 (rst, clk, r23_out, r24_out);
	reg32 r25 (rst, clk, r24_out, r25_out);
	reg32 r26 (rst, clk, r25_out, r26_out);
	reg32 r27 (rst, clk, r26_out, r27_out);
	reg32 r28 (rst, clk, r27_out, r28_out);
	reg32 r29 (rst, clk, r28_out, r29_out);
	reg32 r30 (rst, clk, r29_out, r30_out);
	reg32 r31 (rst, clk, r30_out, r31_out);
	reg32 r32 (rst, clk, r31_out, r32_out);
	reg32 r33 (rst, clk, r32_out, r33_out);
	reg32 r34 (rst, clk, r33_out, r34_out);
	reg32 r35 (rst, clk, r34_out, r35_out);
	reg32 r36 (rst, clk, r35_out, r36_out);
	reg32 r37 (rst, clk, r36_out, r37_out);
	reg32 r38 (rst, clk, r37_out, r38_out);
	reg32 r39 (rst, clk, r38_out, r39_out);
	reg32 r40 (rst, clk, r39_out, r40_out);
	reg32 r41 (rst, clk, r40_out, r41_out);
	reg32 r42 (rst, clk, r41_out, r42_out);
	reg32 r43 (rst, clk, r42_out, r43_out);
	reg32 r44 (rst, clk, r43_out, r44_out);
	reg32 r45 (rst, clk, r44_out, r45_out);
	reg32 r46 (rst, clk, r45_out, r46_out);
	reg32 r47 (rst, clk, r46_out, r47_out);
	reg32 r48 (rst, clk, r47_out, r48_out);
	reg32 r49 (rst, clk, r48_out, r49_out);
	reg32 r50 (rst, clk, r49_out, r50_out);
	reg32 r51 (rst, clk, r50_out, r51_out);
	reg32 r52 (rst, clk, r51_out, r52_out);
	reg32 r53 (rst, clk, r52_out, r53_out);
	reg32 r54 (rst, clk, r53_out, r54_out);
	reg32 r55 (rst, clk, r54_out, r55_out);
	reg32 r56 (rst, clk, r55_out, r56_out);
	reg32 r57 (rst, clk, r56_out, r57_out);
	reg32 r58 (rst, clk, r57_out, r58_out);
	reg32 r59 (rst, clk, r58_out, r59_out);
	reg32 r60 (rst, clk, r59_out, r60_out);
	reg32 r61 (rst, clk, r60_out, r61_out);
	reg32 r62 (rst, clk, r61_out, r62_out);
	reg32 r63 (rst, clk, r62_out, r63_out);
	reg32 r64 (rst, clk, r63_out, r64_out);
	reg32 r65 (rst, clk, r64_out, r65_out);
	reg32 r66 (rst, clk, r65_out, r66_out);
	reg32 r67 (rst, clk, r66_out, r67_out);
	reg32 r68 (rst, clk, r67_out, r68_out);
	reg32 r69 (rst, clk, r68_out, r69_out);
	reg32 r70 (rst, clk, r69_out, r70_out);
	reg32 r71 (rst, clk, r70_out, r71_out);
	reg32 r72 (rst, clk, r71_out, r72_out);
	reg32 r73 (rst, clk, r72_out, r73_out);
	reg32 r74 (rst, clk, r73_out, r74_out);
	reg32 r75 (rst, clk, r74_out, r75_out);
	reg32 r76 (rst, clk, r75_out, r76_out);
	reg32 r77 (rst, clk, r76_out, r77_out);
	reg32 r78 (rst, clk, r77_out, r78_out);
	reg32 r79 (rst, clk, r78_out, r79_out);
	reg32 r80 (rst, clk, r79_out, r80_out);
	reg32 r81 (rst, clk, r80_out, r81_out);
	reg32 r82 (rst, clk, r81_out, r82_out);
	reg32 r83 (rst, clk, r82_out, r83_out);
	reg32 r84 (rst, clk, r83_out, r84_out);
	reg32 r85 (rst, clk, r84_out, r85_out);
	reg32 r86 (rst, clk, r85_out, r86_out);
	reg32 r87 (rst, clk, r86_out, r87_out);
	reg32 r88 (rst, clk, r87_out, r88_out);
	reg32 r89 (rst, clk, r88_out, r89_out);
	reg32 r90 (rst, clk, r89_out, r90_out);
	reg32 r91 (rst, clk, r90_out, r91_out);
	reg32 r92 (rst, clk, r91_out, r92_out);
	reg32 r93 (rst, clk, r92_out, r93_out);
	reg32 r94 (rst, clk, r93_out, r94_out);
	reg32 r95 (rst, clk, r94_out, r95_out);
	reg32 r96 (rst, clk, r95_out, r96_out);
	reg32 r97 (rst, clk, r96_out, r97_out);
	reg32 r98 (rst, clk, r97_out, r98_out);
	reg32 r99 (rst, clk, r98_out, r99_out);
	reg32 r100 (rst, clk, r99_out, r100_out);
	reg32 r101 (rst, clk, r100_out, r101_out);
	reg32 r102 (rst, clk, r101_out, r102_out);
	reg32 r103 (rst, clk, r102_out, r103_out);
	reg32 r104 (rst, clk, r103_out, r104_out);
	reg32 r105 (rst, clk, r104_out, r105_out);
	reg32 r106 (rst, clk, r105_out, r106_out);
	reg32 r107 (rst, clk, r106_out, r107_out);
	reg32 r108 (rst, clk, r107_out, r108_out);
	reg32 r109 (rst, clk, r108_out, r109_out);
	reg32 r110 (rst, clk, r109_out, r110_out);
	reg32 r111 (rst, clk, r110_out, r111_out);
	reg32 r112 (rst, clk, r111_out, r112_out);
	reg32 r113 (rst, clk, r112_out, r113_out);
	reg32 r114 (rst, clk, r113_out, r114_out);
	reg32 r115 (rst, clk, r114_out, r115_out);
	reg32 r116 (rst, clk, r115_out, r116_out);
	reg32 r117 (rst, clk, r116_out, r117_out);
	reg32 r118 (rst, clk, r117_out, r118_out);
	reg32 r119 (rst, clk, r118_out, r119_out);
	reg32 r120 (rst, clk, r119_out, r120_out);
	reg32 r121 (rst, clk, r120_out, r121_out);
	reg32 r122 (rst, clk, r121_out, r122_out);
	reg32 r123 (rst, clk, r122_out, r123_out);
	reg32 r124 (rst, clk, r123_out, r124_out);
	reg32 r125 (rst, clk, r124_out, r125_out);
	reg32 r126 (rst, clk, r125_out, r126_out);
	reg32 r127 (rst, clk, r126_out, r127_out);
	reg32 r128 (rst, clk, r127_out, r128_out);
	reg32 r129 (rst, clk, r128_out, r129_out);
	reg32 r130 (rst, clk, r129_out, r130_out);
	reg32 r131 (rst, clk, r130_out, r131_out);
	reg32 r132 (rst, clk, r131_out, r132_out);
	reg32 r133 (rst, clk, r132_out, r133_out);
	reg32 r134 (rst, clk, r133_out, r134_out);
	reg32 r135 (rst, clk, r134_out, r135_out);
	reg32 r136 (rst, clk, r135_out, r136_out);
	reg32 r137 (rst, clk, r136_out, r137_out);
	reg32 r138 (rst, clk, r137_out, r138_out);
	reg32 r139 (rst, clk, r138_out, r139_out);
	reg32 r140 (rst, clk, r139_out, r140_out);
	reg32 r141 (rst, clk, r140_out, r141_out);
	reg32 r142 (rst, clk, r141_out, r142_out);
	reg32 r143 (rst, clk, r142_out, r143_out);
	reg32 r144 (rst, clk, r143_out, r144_out);
	reg32 r145 (rst, clk, r144_out, r145_out);
	reg32 r146 (rst, clk, r145_out, r146_out);
	reg32 r147 (rst, clk, r146_out, r147_out);
	reg32 r148 (rst, clk, r147_out, r148_out);
	reg32 r149 (rst, clk, r148_out, r149_out);
	reg32 r150 (rst, clk, r149_out, r150_out);
	reg32 r151 (rst, clk, r150_out, r151_out);
	reg32 r152 (rst, clk, r151_out, r152_out);
	reg32 r153 (rst, clk, r152_out, r153_out);
	reg32 r154 (rst, clk, r153_out, r154_out);
	reg32 r155 (rst, clk, r154_out, r155_out);
	reg32 r156 (rst, clk, r155_out, r156_out);
	reg32 r157 (rst, clk, r156_out, r157_out);
	reg32 r158 (rst, clk, r157_out, r158_out);
	reg32 r159 (rst, clk, r158_out, r159_out);
	reg32 r160 (rst, clk, r159_out, r160_out);
	reg32 r161 (rst, clk, r160_out, r161_out);
	reg32 r162 (rst, clk, r161_out, r162_out);
	reg32 r163 (rst, clk, r162_out, r163_out);
	reg32 r164 (rst, clk, r163_out, r164_out);
	reg32 r165 (rst, clk, r164_out, r165_out);
	reg32 r166 (rst, clk, r165_out, r166_out);
	reg32 r167 (rst, clk, r166_out, r167_out);
	reg32 r168 (rst, clk, r167_out, r168_out);
	reg32 r169 (rst, clk, r168_out, r169_out);
	reg32 r170 (rst, clk, r169_out, r170_out);
	reg32 r171 (rst, clk, r170_out, r171_out);
	reg32 r172 (rst, clk, r171_out, r172_out);
	reg32 r173 (rst, clk, r172_out, r173_out);
	reg32 r174 (rst, clk, r173_out, r174_out);
	reg32 r175 (rst, clk, r174_out, r175_out);
	reg32 r176 (rst, clk, r175_out, r176_out);
	reg32 r177 (rst, clk, r176_out, r177_out);
	reg32 r178 (rst, clk, r177_out, r178_out);
	reg32 r179 (rst, clk, r178_out, r179_out);
	reg32 r180 (rst, clk, r179_out, r180_out);
	reg32 r181 (rst, clk, r180_out, r181_out);
	reg32 r182 (rst, clk, r181_out, r182_out);
	reg32 r183 (rst, clk, r182_out, r183_out);
	reg32 r184 (rst, clk, r183_out, r184_out);
	reg32 r185 (rst, clk, r184_out, r185_out);
	reg32 r186 (rst, clk, r185_out, r186_out);
	reg32 r187 (rst, clk, r186_out, r187_out);
	reg32 r188 (rst, clk, r187_out, r188_out);
	reg32 r189 (rst, clk, r188_out, r189_out);
	reg32 r190 (rst, clk, r189_out, r190_out);
	reg32 r191 (rst, clk, r190_out, r191_out);
	reg32 r192 (rst, clk, r191_out, r192_out);
	reg32 r193 (rst, clk, r192_out, r193_out);
	reg32 r194 (rst, clk, r193_out, r194_out);
	reg32 r195 (rst, clk, r194_out, r195_out);
	reg32 r196 (rst, clk, r195_out, r196_out);
	reg32 r197 (rst, clk, r196_out, r197_out);
	reg32 r198 (rst, clk, r197_out, r198_out);
	reg32 r199 (rst, clk, r198_out, r199_out);
	reg32 r200 (rst, clk, r199_out, r200_out);
	reg32 r201 (rst, clk, r200_out, r201_out);
	reg32 r202 (rst, clk, r201_out, r202_out);
	reg32 r203 (rst, clk, r202_out, r203_out);
	reg32 r204 (rst, clk, r203_out, r204_out);
	reg32 r205 (rst, clk, r204_out, r205_out);
	reg32 r206 (rst, clk, r205_out, r206_out);
	reg32 r207 (rst, clk, r206_out, r207_out);
	reg32 r208 (rst, clk, r207_out, r208_out);
	reg32 r209 (rst, clk, r208_out, r209_out);
	reg32 r210 (rst, clk, r209_out, r210_out);
	reg32 r211 (rst, clk, r210_out, r211_out);
	reg32 r212 (rst, clk, r211_out, r212_out);
	reg32 r213 (rst, clk, r212_out, r213_out);
	reg32 r214 (rst, clk, r213_out, r214_out);
	reg32 r215 (rst, clk, r214_out, r215_out);
	reg32 r216 (rst, clk, r215_out, r216_out);
	reg32 r217 (rst, clk, r216_out, r217_out);
	reg32 r218 (rst, clk, r217_out, r218_out);
	reg32 r219 (rst, clk, r218_out, r219_out);
	reg32 r220 (rst, clk, r219_out, r220_out);
	reg32 r221 (rst, clk, r220_out, r221_out);
	reg32 r222 (rst, clk, r221_out, r222_out);
	reg32 r223 (rst, clk, r222_out, r223_out);
	reg32 r224 (rst, clk, r223_out, r224_out);
	reg32 r225 (rst, clk, r224_out, r225_out);
	reg32 r226 (rst, clk, r225_out, r226_out);
	reg32 r227 (rst, clk, r226_out, r227_out);
	reg32 r228 (rst, clk, r227_out, r228_out);
	reg32 r229 (rst, clk, r228_out, r229_out);
	reg32 r230 (rst, clk, r229_out, r230_out);
	reg32 r231 (rst, clk, r230_out, r231_out);
	reg32 r232 (rst, clk, r231_out, r232_out);
	reg32 r233 (rst, clk, r232_out, r233_out);
	reg32 r234 (rst, clk, r233_out, r234_out);
	reg32 r235 (rst, clk, r234_out, r235_out);
	reg32 r236 (rst, clk, r235_out, r236_out);
	reg32 r237 (rst, clk, r236_out, r237_out);
	reg32 r238 (rst, clk, r237_out, r238_out);
	reg32 r239 (rst, clk, r238_out, r239_out);
	reg32 r240 (rst, clk, r239_out, r240_out);
	reg32 r241 (rst, clk, r240_out, r241_out);
	reg32 r242 (rst, clk, r241_out, r242_out);
	reg32 r243 (rst, clk, r242_out, r243_out);
	reg32 r244 (rst, clk, r243_out, r244_out);
	reg32 r245 (rst, clk, r244_out, r245_out);
	reg32 r246 (rst, clk, r245_out, r246_out);
	reg32 r247 (rst, clk, r246_out, r247_out);
	reg32 r248 (rst, clk, r247_out, r248_out);
	reg32 r249 (rst, clk, r248_out, r249_out);
	reg32 r250 (rst, clk, r249_out, r250_out);
	reg32 r251 (rst, clk, r250_out, r251_out);
	reg32 r252 (rst, clk, r251_out, r252_out);
	reg32 r253 (rst, clk, r252_out, r253_out);
	reg32 r254 (rst, clk, r253_out, r254_out);
	reg32 r255 (rst, clk, r254_out, r255_out);
	reg32 r256 (rst, clk, r255_out, r256_out);
	reg32 r257 (rst, clk, r256_out, r257_out);
	reg32 r258 (rst, clk, r257_out, r258_out);
	reg32 r259 (rst, clk, r258_out, r259_out);
	reg32 r260 (rst, clk, r259_out, r260_out);
	reg32 r261 (rst, clk, r260_out, r261_out);
	reg32 r262 (rst, clk, r261_out, r262_out);
	reg32 r263 (rst, clk, r262_out, r263_out);
	reg32 r264 (rst, clk, r263_out, r264_out);
	reg32 r265 (rst, clk, r264_out, r265_out);
	reg32 r266 (rst, clk, r265_out, r266_out);
	reg32 r267 (rst, clk, r266_out, r267_out);
	reg32 r268 (rst, clk, r267_out, r268_out);
	reg32 r269 (rst, clk, r268_out, r269_out);
	reg32 r270 (rst, clk, r269_out, r270_out);
	reg32 r271 (rst, clk, r270_out, r271_out);
	reg32 r272 (rst, clk, r271_out, r272_out);
	reg32 r273 (rst, clk, r272_out, r273_out);
	reg32 r274 (rst, clk, r273_out, r274_out);
	reg32 r275 (rst, clk, r274_out, r275_out);
	reg32 r276 (rst, clk, r275_out, r276_out);
	reg32 r277 (rst, clk, r276_out, r277_out);
	reg32 r278 (rst, clk, r277_out, r278_out);
	reg32 r279 (rst, clk, r278_out, r279_out);
	reg32 r280 (rst, clk, r279_out, r280_out);
	reg32 r281 (rst, clk, r280_out, r281_out);
	reg32 r282 (rst, clk, r281_out, r282_out);
	reg32 r283 (rst, clk, r282_out, r283_out);
	reg32 r284 (rst, clk, r283_out, r284_out);
	reg32 r285 (rst, clk, r284_out, r285_out);
	reg32 r286 (rst, clk, r285_out, r286_out);
	reg32 r287 (rst, clk, r286_out, r287_out);
	reg32 r288 (rst, clk, r287_out, r288_out);
	reg32 r289 (rst, clk, r288_out, r289_out);
	reg32 r290 (rst, clk, r289_out, r290_out);
	reg32 r291 (rst, clk, r290_out, r291_out);
	reg32 r292 (rst, clk, r291_out, r292_out);
	reg32 r293 (rst, clk, r292_out, r293_out);
	reg32 r294 (rst, clk, r293_out, r294_out);
	reg32 r295 (rst, clk, r294_out, r295_out);
	reg32 r296 (rst, clk, r295_out, r296_out);
	reg32 r297 (rst, clk, r296_out, r297_out);
	reg32 r298 (rst, clk, r297_out, r298_out);
	reg32 r299 (rst, clk, r298_out, r299_out);
	reg32 r300 (rst, clk, r299_out, r300_out);
	reg32 r301 (rst, clk, r300_out, r301_out);
	reg32 r302 (rst, clk, r301_out, r302_out);
	reg32 r303 (rst, clk, r302_out, r303_out);
	reg32 r304 (rst, clk, r303_out, r304_out);
	reg32 r305 (rst, clk, r304_out, r305_out);
	reg32 r306 (rst, clk, r305_out, r306_out);
	reg32 r307 (rst, clk, r306_out, r307_out);
	reg32 r308 (rst, clk, r307_out, r308_out);
	reg32 r309 (rst, clk, r308_out, r309_out);
	reg32 r310 (rst, clk, r309_out, r310_out);
	reg32 r311 (rst, clk, r310_out, r311_out);
	reg32 r312 (rst, clk, r311_out, r312_out);
	reg32 r313 (rst, clk, r312_out, r313_out);
	reg32 r314 (rst, clk, r313_out, r314_out);
	reg32 r315 (rst, clk, r314_out, r315_out);
	reg32 r316 (rst, clk, r315_out, r316_out);
	reg32 r317 (rst, clk, r316_out, r317_out);
	reg32 r318 (rst, clk, r317_out, r318_out);
	reg32 r319 (rst, clk, r318_out, r319_out);
	reg32 r320 (rst, clk, r319_out, r320_out);
	reg32 r321 (rst, clk, r320_out, r321_out);
	reg32 r322 (rst, clk, r321_out, r322_out);
	reg32 r323 (rst, clk, r322_out, r323_out);
	reg32 r324 (rst, clk, r323_out, r324_out);
	reg32 r325 (rst, clk, r324_out, r325_out);
	reg32 r326 (rst, clk, r325_out, r326_out);
	reg32 r327 (rst, clk, r326_out, r327_out);
	reg32 r328 (rst, clk, r327_out, r328_out);
	reg32 r329 (rst, clk, r328_out, r329_out);
	reg32 r330 (rst, clk, r329_out, r330_out);
	reg32 r331 (rst, clk, r330_out, r331_out);
	reg32 r332 (rst, clk, r331_out, r332_out);
	reg32 r333 (rst, clk, r332_out, r333_out);
	reg32 r334 (rst, clk, r333_out, r334_out);
	reg32 r335 (rst, clk, r334_out, r335_out);
	reg32 r336 (rst, clk, r335_out, r336_out);
	reg32 r337 (rst, clk, r336_out, r337_out);
	reg32 r338 (rst, clk, r337_out, r338_out);
	reg32 r339 (rst, clk, r338_out, r339_out);
	reg32 r340 (rst, clk, r339_out, r340_out);
	reg32 r341 (rst, clk, r340_out, r341_out);
	reg32 r342 (rst, clk, r341_out, r342_out);
	reg32 r343 (rst, clk, r342_out, r343_out);
	reg32 r344 (rst, clk, r343_out, r344_out);
	reg32 r345 (rst, clk, r344_out, r345_out);
	reg32 r346 (rst, clk, r345_out, r346_out);
	reg32 r347 (rst, clk, r346_out, r347_out);
	reg32 r348 (rst, clk, r347_out, r348_out);
	reg32 r349 (rst, clk, r348_out, r349_out);
	reg32 r350 (rst, clk, r349_out, r350_out);
	reg32 r351 (rst, clk, r350_out, r351_out);
	reg32 r352 (rst, clk, r351_out, r352_out);
	reg32 r353 (rst, clk, r352_out, r353_out);
	reg32 r354 (rst, clk, r353_out, r354_out);
	reg32 r355 (rst, clk, r354_out, r355_out);
	reg32 r356 (rst, clk, r355_out, r356_out);
	reg32 r357 (rst, clk, r356_out, r357_out);
	reg32 r358 (rst, clk, r357_out, r358_out);
	reg32 r359 (rst, clk, r358_out, r359_out);
	reg32 r360 (rst, clk, r359_out, r360_out);
	reg32 r361 (rst, clk, r360_out, r361_out);
	reg32 r362 (rst, clk, r361_out, r362_out);
	reg32 r363 (rst, clk, r362_out, r363_out);
	reg32 r364 (rst, clk, r363_out, r364_out);
	reg32 r365 (rst, clk, r364_out, r365_out);
	reg32 r366 (rst, clk, r365_out, r366_out);
	reg32 r367 (rst, clk, r366_out, r367_out);
	reg32 r368 (rst, clk, r367_out, r368_out);
	reg32 r369 (rst, clk, r368_out, r369_out);
	reg32 r370 (rst, clk, r369_out, r370_out);
	reg32 r371 (rst, clk, r370_out, r371_out);
	reg32 r372 (rst, clk, r371_out, r372_out);
	reg32 r373 (rst, clk, r372_out, r373_out);
	reg32 r374 (rst, clk, r373_out, r374_out);
	reg32 r375 (rst, clk, r374_out, r375_out);
	reg32 r376 (rst, clk, r375_out, r376_out);
	reg32 r377 (rst, clk, r376_out, r377_out);
	reg32 r378 (rst, clk, r377_out, r378_out);
	reg32 r379 (rst, clk, r378_out, r379_out);
	reg32 r380 (rst, clk, r379_out, r380_out);
	reg32 r381 (rst, clk, r380_out, r381_out);
	reg32 r382 (rst, clk, r381_out, r382_out);
	reg32 r383 (rst, clk, r382_out, r383_out);
	reg32 r384 (rst, clk, r383_out, r384_out);
	reg32 r385 (rst, clk, r384_out, r385_out);
	reg32 r386 (rst, clk, r385_out, r386_out);
	reg32 r387 (rst, clk, r386_out, r387_out);
	reg32 r388 (rst, clk, r387_out, r388_out);
	reg32 r389 (rst, clk, r388_out, r389_out);
	reg32 r390 (rst, clk, r389_out, r390_out);
	reg32 r391 (rst, clk, r390_out, r391_out);
	reg32 r392 (rst, clk, r391_out, r392_out);
	reg32 r393 (rst, clk, r392_out, r393_out);
	reg32 r394 (rst, clk, r393_out, r394_out);
	reg32 r395 (rst, clk, r394_out, r395_out);
	reg32 r396 (rst, clk, r395_out, r396_out);
	reg32 r397 (rst, clk, r396_out, r397_out);
	reg32 r398 (rst, clk, r397_out, r398_out);
	reg32 r399 (rst, clk, r398_out, r399_out);
	reg32 r400 (rst, clk, r399_out, r400_out);
	reg32 r401 (rst, clk, r400_out, r401_out);
	reg32 r402 (rst, clk, r401_out, r402_out);
	reg32 r403 (rst, clk, r402_out, r403_out);
	reg32 r404 (rst, clk, r403_out, r404_out);
	reg32 r405 (rst, clk, r404_out, r405_out);
	reg32 r406 (rst, clk, r405_out, r406_out);
	reg32 r407 (rst, clk, r406_out, r407_out);
	reg32 r408 (rst, clk, r407_out, r408_out);
	reg32 r409 (rst, clk, r408_out, r409_out);
	reg32 r410 (rst, clk, r409_out, r410_out);
	reg32 r411 (rst, clk, r410_out, r411_out);
	reg32 r412 (rst, clk, r411_out, r412_out);
	reg32 r413 (rst, clk, r412_out, r413_out);
	reg32 r414 (rst, clk, r413_out, r414_out);
	reg32 r415 (rst, clk, r414_out, r415_out);
	reg32 r416 (rst, clk, r415_out, r416_out);
	reg32 r417 (rst, clk, r416_out, r417_out);
	reg32 r418 (rst, clk, r417_out, r418_out);
	reg32 r419 (rst, clk, r418_out, r419_out);
	reg32 r420 (rst, clk, r419_out, r420_out);
	reg32 r421 (rst, clk, r420_out, r421_out);
	reg32 r422 (rst, clk, r421_out, r422_out);
	reg32 r423 (rst, clk, r422_out, r423_out);
	reg32 r424 (rst, clk, r423_out, r424_out);
	reg32 r425 (rst, clk, r424_out, r425_out);
	reg32 r426 (rst, clk, r425_out, r426_out);
	reg32 r427 (rst, clk, r426_out, r427_out);
	reg32 r428 (rst, clk, r427_out, r428_out);
	reg32 r429 (rst, clk, r428_out, r429_out);
	reg32 r430 (rst, clk, r429_out, r430_out);
	reg32 r431 (rst, clk, r430_out, r431_out);
	reg32 r432 (rst, clk, r431_out, r432_out);
	reg32 r433 (rst, clk, r432_out, r433_out);
	reg32 r434 (rst, clk, r433_out, r434_out);
	reg32 r435 (rst, clk, r434_out, r435_out);
	reg32 r436 (rst, clk, r435_out, r436_out);
	reg32 r437 (rst, clk, r436_out, r437_out);
	reg32 r438 (rst, clk, r437_out, r438_out);
	reg32 r439 (rst, clk, r438_out, r439_out);
	reg32 r440 (rst, clk, r439_out, r440_out);
	reg32 r441 (rst, clk, r440_out, r441_out);
	reg32 r442 (rst, clk, r441_out, r442_out);
	reg32 r443 (rst, clk, r442_out, r443_out);
	reg32 r444 (rst, clk, r443_out, r444_out);
	reg32 r445 (rst, clk, r444_out, r445_out);
	reg32 r446 (rst, clk, r445_out, r446_out);
	reg32 r447 (rst, clk, r446_out, r447_out);
	reg32 r448 (rst, clk, r447_out, r448_out);
	reg32 r449 (rst, clk, r448_out, r449_out);
	reg32 r450 (rst, clk, r449_out, r450_out);
	reg32 r451 (rst, clk, r450_out, r451_out);
	reg32 r452 (rst, clk, r451_out, r452_out);
	reg32 r453 (rst, clk, r452_out, r453_out);
	reg32 r454 (rst, clk, r453_out, r454_out);
	reg32 r455 (rst, clk, r454_out, r455_out);
	reg32 r456 (rst, clk, r455_out, r456_out);
	reg32 r457 (rst, clk, r456_out, r457_out);
	reg32 r458 (rst, clk, r457_out, r458_out);
	reg32 r459 (rst, clk, r458_out, r459_out);
	reg32 r460 (rst, clk, r459_out, r460_out);
	reg32 r461 (rst, clk, r460_out, r461_out);
	reg32 r462 (rst, clk, r461_out, r462_out);
	reg32 r463 (rst, clk, r462_out, r463_out);
	reg32 r464 (rst, clk, r463_out, r464_out);
	reg32 r465 (rst, clk, r464_out, r465_out);
	reg32 r466 (rst, clk, r465_out, r466_out);
	reg32 r467 (rst, clk, r466_out, r467_out);
	reg32 r468 (rst, clk, r467_out, r468_out);
	reg32 r469 (rst, clk, r468_out, r469_out);
	reg32 r470 (rst, clk, r469_out, r470_out);
	reg32 r471 (rst, clk, r470_out, r471_out);
	reg32 r472 (rst, clk, r471_out, r472_out);
	reg32 r473 (rst, clk, r472_out, r473_out);
	reg32 r474 (rst, clk, r473_out, r474_out);
	reg32 r475 (rst, clk, r474_out, r475_out);
	reg32 r476 (rst, clk, r475_out, r476_out);
	reg32 r477 (rst, clk, r476_out, r477_out);
	reg32 r478 (rst, clk, r477_out, r478_out);
	reg32 r479 (rst, clk, r478_out, r479_out);
	reg32 r480 (rst, clk, r479_out, r480_out);
	reg32 r481 (rst, clk, r480_out, r481_out);
	reg32 r482 (rst, clk, r481_out, r482_out);
	reg32 r483 (rst, clk, r482_out, r483_out);
	reg32 r484 (rst, clk, r483_out, r484_out);
	reg32 r485 (rst, clk, r484_out, r485_out);
	reg32 r486 (rst, clk, r485_out, r486_out);
	reg32 r487 (rst, clk, r486_out, r487_out);
	reg32 r488 (rst, clk, r487_out, r488_out);
	reg32 r489 (rst, clk, r488_out, r489_out);
	reg32 r490 (rst, clk, r489_out, r490_out);
	reg32 r491 (rst, clk, r490_out, r491_out);
	reg32 r492 (rst, clk, r491_out, r492_out);
	reg32 r493 (rst, clk, r492_out, r493_out);
	reg32 r494 (rst, clk, r493_out, r494_out);
	reg32 r495 (rst, clk, r494_out, r495_out);
	reg32 r496 (rst, clk, r495_out, r496_out);
	reg32 r497 (rst, clk, r496_out, r497_out);
	reg32 r498 (rst, clk, r497_out, r498_out);
	reg32 r499 (rst, clk, r498_out, r499_out);
	reg32 r500 (rst, clk, r499_out, r500_out);
	reg32 r501 (rst, clk, r500_out, r501_out);
	reg32 r502 (rst, clk, r501_out, r502_out);
	reg32 r503 (rst, clk, r502_out, r503_out);
	reg32 r504 (rst, clk, r503_out, r504_out);
	reg32 r505 (rst, clk, r504_out, r505_out);
	reg32 r506 (rst, clk, r505_out, r506_out);
	reg32 r507 (rst, clk, r506_out, r507_out);
	reg32 r508 (rst, clk, r507_out, r508_out);
	reg32 r509 (rst, clk, r508_out, r509_out);
	reg32 r510 (rst, clk, r509_out, r510_out);
	reg32 r511 (rst, clk, r510_out, r511_out);
	reg32 r512 (rst, clk, r511_out, r512_out);
	reg32 r513 (rst, clk, r512_out, r513_out);
	reg32 r514 (rst, clk, r513_out, r514_out);
	reg32 r515 (rst, clk, r514_out, r515_out);
	reg32 r516 (rst, clk, r515_out, r516_out);
	reg32 r517 (rst, clk, r516_out, r517_out);
	reg32 r518 (rst, clk, r517_out, r518_out);
	reg32 r519 (rst, clk, r518_out, r519_out);
	reg32 r520 (rst, clk, r519_out, r520_out);
	reg32 r521 (rst, clk, r520_out, r521_out);
	reg32 r522 (rst, clk, r521_out, r522_out);
	reg32 r523 (rst, clk, r522_out, r523_out);
	reg32 r524 (rst, clk, r523_out, r524_out);
	reg32 r525 (rst, clk, r524_out, r525_out);
	reg32 r526 (rst, clk, r525_out, r526_out);
	reg32 r527 (rst, clk, r526_out, r527_out);
	reg32 r528 (rst, clk, r527_out, r528_out);
	reg32 r529 (rst, clk, r528_out, r529_out);
	reg32 r530 (rst, clk, r529_out, r530_out);
	reg32 r531 (rst, clk, r530_out, r531_out);
	reg32 r532 (rst, clk, r531_out, r532_out);
	reg32 r533 (rst, clk, r532_out, r533_out);
	reg32 r534 (rst, clk, r533_out, r534_out);
	reg32 r535 (rst, clk, r534_out, r535_out);
	reg32 r536 (rst, clk, r535_out, r536_out);
	reg32 r537 (rst, clk, r536_out, r537_out);
	reg32 r538 (rst, clk, r537_out, r538_out);
	reg32 r539 (rst, clk, r538_out, r539_out);
	reg32 r540 (rst, clk, r539_out, r540_out);
	reg32 r541 (rst, clk, r540_out, r541_out);
	reg32 r542 (rst, clk, r541_out, r542_out);
	reg32 r543 (rst, clk, r542_out, r543_out);
	reg32 r544 (rst, clk, r543_out, r544_out);
	reg32 r545 (rst, clk, r544_out, r545_out);
	reg32 r546 (rst, clk, r545_out, r546_out);
	reg32 r547 (rst, clk, r546_out, r547_out);
	reg32 r548 (rst, clk, r547_out, r548_out);
	reg32 r549 (rst, clk, r548_out, r549_out);
	reg32 r550 (rst, clk, r549_out, r550_out);
	reg32 r551 (rst, clk, r550_out, r551_out);
	reg32 r552 (rst, clk, r551_out, r552_out);
	reg32 r553 (rst, clk, r552_out, r553_out);
	reg32 r554 (rst, clk, r553_out, r554_out);
	reg32 r555 (rst, clk, r554_out, r555_out);
	reg32 r556 (rst, clk, r555_out, r556_out);
	reg32 r557 (rst, clk, r556_out, r557_out);
	reg32 r558 (rst, clk, r557_out, r558_out);
	reg32 r559 (rst, clk, r558_out, r559_out);
	reg32 r560 (rst, clk, r559_out, r560_out);
	reg32 r561 (rst, clk, r560_out, r561_out);
	reg32 r562 (rst, clk, r561_out, r562_out);
	reg32 r563 (rst, clk, r562_out, r563_out);
	reg32 r564 (rst, clk, r563_out, r564_out);
	reg32 r565 (rst, clk, r564_out, r565_out);
	reg32 r566 (rst, clk, r565_out, r566_out);
	reg32 r567 (rst, clk, r566_out, r567_out);
	reg32 r568 (rst, clk, r567_out, r568_out);
	reg32 r569 (rst, clk, r568_out, r569_out);
	reg32 r570 (rst, clk, r569_out, r570_out);
	reg32 r571 (rst, clk, r570_out, r571_out);
	reg32 r572 (rst, clk, r571_out, r572_out);
	reg32 r573 (rst, clk, r572_out, r573_out);
	reg32 r574 (rst, clk, r573_out, r574_out);
	reg32 r575 (rst, clk, r574_out, r575_out);
	reg32 r576 (rst, clk, r575_out, r576_out);
	reg32 r577 (rst, clk, r576_out, r577_out);
	reg32 r578 (rst, clk, r577_out, r578_out);
	reg32 r579 (rst, clk, r578_out, r579_out);
	reg32 r580 (rst, clk, r579_out, r580_out);
	reg32 r581 (rst, clk, r580_out, r581_out);
	reg32 r582 (rst, clk, r581_out, r582_out);
	reg32 r583 (rst, clk, r582_out, r583_out);
	reg32 r584 (rst, clk, r583_out, r584_out);
	reg32 r585 (rst, clk, r584_out, r585_out);
	reg32 r586 (rst, clk, r585_out, r586_out);
	reg32 r587 (rst, clk, r586_out, r587_out);
	reg32 r588 (rst, clk, r587_out, r588_out);
	reg32 r589 (rst, clk, r588_out, r589_out);
	reg32 r590 (rst, clk, r589_out, r590_out);
	reg32 r591 (rst, clk, r590_out, r591_out);
	reg32 r592 (rst, clk, r591_out, r592_out);
	reg32 r593 (rst, clk, r592_out, r593_out);
	reg32 r594 (rst, clk, r593_out, r594_out);
	reg32 r595 (rst, clk, r594_out, r595_out);
	reg32 r596 (rst, clk, r595_out, r596_out);
	reg32 r597 (rst, clk, r596_out, r597_out);
	reg32 r598 (rst, clk, r597_out, r598_out);
	reg32 r599 (rst, clk, r598_out, r599_out);
	reg32 r600 (rst, clk, r599_out, r600_out);
	reg32 r601 (rst, clk, r600_out, r601_out);
	reg32 r602 (rst, clk, r601_out, r602_out);
	reg32 r603 (rst, clk, r602_out, r603_out);
	reg32 r604 (rst, clk, r603_out, r604_out);
	reg32 r605 (rst, clk, r604_out, r605_out);
	reg32 r606 (rst, clk, r605_out, r606_out);
	reg32 r607 (rst, clk, r606_out, r607_out);
	reg32 r608 (rst, clk, r607_out, r608_out);
	reg32 r609 (rst, clk, r608_out, r609_out);
	reg32 r610 (rst, clk, r609_out, r610_out);
	reg32 r611 (rst, clk, r610_out, r611_out);
	reg32 r612 (rst, clk, r611_out, r612_out);
	reg32 r613 (rst, clk, r612_out, r613_out);
	reg32 r614 (rst, clk, r613_out, r614_out);
	reg32 r615 (rst, clk, r614_out, r615_out);
	reg32 r616 (rst, clk, r615_out, r616_out);
	reg32 r617 (rst, clk, r616_out, r617_out);
	reg32 r618 (rst, clk, r617_out, r618_out);
	reg32 r619 (rst, clk, r618_out, r619_out);
	reg32 r620 (rst, clk, r619_out, r620_out);
	reg32 r621 (rst, clk, r620_out, r621_out);
	reg32 r622 (rst, clk, r621_out, r622_out);
	reg32 r623 (rst, clk, r622_out, r623_out);
	reg32 r624 (rst, clk, r623_out, r624_out);
	reg32 r625 (rst, clk, r624_out, r625_out);
	reg32 r626 (rst, clk, r625_out, r626_out);
	reg32 r627 (rst, clk, r626_out, r627_out);
	reg32 r628 (rst, clk, r627_out, r628_out);
	reg32 r629 (rst, clk, r628_out, r629_out);
	reg32 r630 (rst, clk, r629_out, r630_out);
	reg32 r631 (rst, clk, r630_out, r631_out);
	reg32 r632 (rst, clk, r631_out, r632_out);
	reg32 r633 (rst, clk, r632_out, r633_out);
	reg32 r634 (rst, clk, r633_out, r634_out);
	reg32 r635 (rst, clk, r634_out, r635_out);
	reg32 r636 (rst, clk, r635_out, r636_out);
	reg32 r637 (rst, clk, r636_out, r637_out);
	reg32 r638 (rst, clk, r637_out, r638_out);
	reg32 r639 (rst, clk, r638_out, r639_out);
	reg32 r640 (rst, clk, r639_out, r640_out);
	reg32 r641 (rst, clk, r640_out, r641_out);
	reg32 r642 (rst, clk, r641_out, r642_out);
	reg32 r643 (rst, clk, r642_out, r643_out);
	reg32 r644 (rst, clk, r643_out, r644_out);
	reg32 r645 (rst, clk, r644_out, r645_out);
	reg32 r646 (rst, clk, r645_out, r646_out);
	reg32 r647 (rst, clk, r646_out, r647_out);
	reg32 r648 (rst, clk, r647_out, r648_out);
	reg32 r649 (rst, clk, r648_out, r649_out);
	reg32 r650 (rst, clk, r649_out, r650_out);
	reg32 r651 (rst, clk, r650_out, r651_out);
	reg32 r652 (rst, clk, r651_out, r652_out);
	reg32 r653 (rst, clk, r652_out, r653_out);
	reg32 r654 (rst, clk, r653_out, r654_out);
	reg32 r655 (rst, clk, r654_out, r655_out);
	reg32 r656 (rst, clk, r655_out, r656_out);
	reg32 r657 (rst, clk, r656_out, r657_out);
	reg32 r658 (rst, clk, r657_out, r658_out);
	reg32 r659 (rst, clk, r658_out, r659_out);
	reg32 r660 (rst, clk, r659_out, r660_out);
	reg32 r661 (rst, clk, r660_out, r661_out);
	reg32 r662 (rst, clk, r661_out, r662_out);
	reg32 r663 (rst, clk, r662_out, r663_out);
	reg32 r664 (rst, clk, r663_out, r664_out);
	reg32 r665 (rst, clk, r664_out, r665_out);
	reg32 r666 (rst, clk, r665_out, r666_out);
	reg32 r667 (rst, clk, r666_out, r667_out);
	reg32 r668 (rst, clk, r667_out, r668_out);
	reg32 r669 (rst, clk, r668_out, r669_out);
	reg32 r670 (rst, clk, r669_out, r670_out);
	reg32 r671 (rst, clk, r670_out, r671_out);
	reg32 r672 (rst, clk, r671_out, r672_out);
	reg32 r673 (rst, clk, r672_out, r673_out);
	reg32 r674 (rst, clk, r673_out, r674_out);
	reg32 r675 (rst, clk, r674_out, r675_out);
	reg32 r676 (rst, clk, r675_out, r676_out);
	reg32 r677 (rst, clk, r676_out, r677_out);
	reg32 r678 (rst, clk, r677_out, r678_out);
	reg32 r679 (rst, clk, r678_out, r679_out);
	reg32 r680 (rst, clk, r679_out, r680_out);
	reg32 r681 (rst, clk, r680_out, r681_out);
	reg32 r682 (rst, clk, r681_out, r682_out);
	reg32 r683 (rst, clk, r682_out, r683_out);
	reg32 r684 (rst, clk, r683_out, r684_out);
	reg32 r685 (rst, clk, r684_out, r685_out);
	reg32 r686 (rst, clk, r685_out, r686_out);
	reg32 r687 (rst, clk, r686_out, r687_out);
	reg32 r688 (rst, clk, r687_out, r688_out);
	reg32 r689 (rst, clk, r688_out, r689_out);
	reg32 r690 (rst, clk, r689_out, r690_out);
	reg32 r691 (rst, clk, r690_out, r691_out);
	reg32 r692 (rst, clk, r691_out, r692_out);
	reg32 r693 (rst, clk, r692_out, r693_out);
	reg32 r694 (rst, clk, r693_out, r694_out);
	reg32 r695 (rst, clk, r694_out, r695_out);
	reg32 r696 (rst, clk, r695_out, r696_out);
	reg32 r697 (rst, clk, r696_out, r697_out);
	reg32 r698 (rst, clk, r697_out, r698_out);
	reg32 r699 (rst, clk, r698_out, r699_out);
	reg32 r700 (rst, clk, r699_out, r700_out);
	reg32 r701 (rst, clk, r700_out, r701_out);
	reg32 r702 (rst, clk, r701_out, r702_out);
	reg32 r703 (rst, clk, r702_out, r703_out);
	reg32 r704 (rst, clk, r703_out, r704_out);
	reg32 r705 (rst, clk, r704_out, r705_out);
	reg32 r706 (rst, clk, r705_out, r706_out);
	reg32 r707 (rst, clk, r706_out, r707_out);
	reg32 r708 (rst, clk, r707_out, r708_out);
	reg32 r709 (rst, clk, r708_out, r709_out);
	reg32 r710 (rst, clk, r709_out, r710_out);
	reg32 r711 (rst, clk, r710_out, r711_out);
	reg32 r712 (rst, clk, r711_out, r712_out);
	reg32 r713 (rst, clk, r712_out, r713_out);
	reg32 r714 (rst, clk, r713_out, r714_out);
	reg32 r715 (rst, clk, r714_out, r715_out);
	reg32 r716 (rst, clk, r715_out, r716_out);
	reg32 r717 (rst, clk, r716_out, r717_out);
	reg32 r718 (rst, clk, r717_out, r718_out);
	reg32 r719 (rst, clk, r718_out, r719_out);
	reg32 r720 (rst, clk, r719_out, r720_out);
	reg32 r721 (rst, clk, r720_out, r721_out);
	reg32 r722 (rst, clk, r721_out, r722_out);
	reg32 r723 (rst, clk, r722_out, r723_out);
	reg32 r724 (rst, clk, r723_out, r724_out);
	reg32 r725 (rst, clk, r724_out, r725_out);
	reg32 r726 (rst, clk, r725_out, r726_out);
	reg32 r727 (rst, clk, r726_out, r727_out);
	reg32 r728 (rst, clk, r727_out, r728_out);
	reg32 r729 (rst, clk, r728_out, r729_out);
	reg32 r730 (rst, clk, r729_out, r730_out);
	reg32 r731 (rst, clk, r730_out, r731_out);
	reg32 r732 (rst, clk, r731_out, r732_out);
	reg32 r733 (rst, clk, r732_out, r733_out);
	reg32 r734 (rst, clk, r733_out, r734_out);
	reg32 r735 (rst, clk, r734_out, r735_out);
	reg32 r736 (rst, clk, r735_out, r736_out);
	reg32 r737 (rst, clk, r736_out, r737_out);
	reg32 r738 (rst, clk, r737_out, r738_out);
	reg32 r739 (rst, clk, r738_out, r739_out);
	reg32 r740 (rst, clk, r739_out, r740_out);
	reg32 r741 (rst, clk, r740_out, r741_out);
	reg32 r742 (rst, clk, r741_out, r742_out);
	reg32 r743 (rst, clk, r742_out, r743_out);
	reg32 r744 (rst, clk, r743_out, r744_out);
	reg32 r745 (rst, clk, r744_out, r745_out);
	reg32 r746 (rst, clk, r745_out, r746_out);
	reg32 r747 (rst, clk, r746_out, r747_out);
	reg32 r748 (rst, clk, r747_out, r748_out);
	reg32 r749 (rst, clk, r748_out, r749_out);
	reg32 r750 (rst, clk, r749_out, r750_out);
	reg32 r751 (rst, clk, r750_out, r751_out);
	reg32 r752 (rst, clk, r751_out, r752_out);
	reg32 r753 (rst, clk, r752_out, r753_out);
	reg32 r754 (rst, clk, r753_out, r754_out);
	reg32 r755 (rst, clk, r754_out, r755_out);
	reg32 r756 (rst, clk, r755_out, r756_out);
	reg32 r757 (rst, clk, r756_out, r757_out);
	reg32 r758 (rst, clk, r757_out, r758_out);
	reg32 r759 (rst, clk, r758_out, r759_out);
	reg32 r760 (rst, clk, r759_out, r760_out);
	reg32 r761 (rst, clk, r760_out, r761_out);
	reg32 r762 (rst, clk, r761_out, r762_out);
	reg32 r763 (rst, clk, r762_out, r763_out);
	reg32 r764 (rst, clk, r763_out, r764_out);
	reg32 r765 (rst, clk, r764_out, r765_out);
	reg32 r766 (rst, clk, r765_out, r766_out);
	reg32 r767 (rst, clk, r766_out, r767_out);
	reg32 r768 (rst, clk, r767_out, r768_out);
	reg32 r769 (rst, clk, r768_out, r769_out);
	reg32 r770 (rst, clk, r769_out, r770_out);
	reg32 r771 (rst, clk, r770_out, r771_out);
	reg32 r772 (rst, clk, r771_out, r772_out);
	reg32 r773 (rst, clk, r772_out, r773_out);
	reg32 r774 (rst, clk, r773_out, r774_out);
	reg32 r775 (rst, clk, r774_out, r775_out);
	reg32 r776 (rst, clk, r775_out, r776_out);
	reg32 r777 (rst, clk, r776_out, r777_out);
	reg32 r778 (rst, clk, r777_out, r778_out);
	reg32 r779 (rst, clk, r778_out, r779_out);
	reg32 r780 (rst, clk, r779_out, r780_out);
	reg32 r781 (rst, clk, r780_out, r781_out);
	reg32 r782 (rst, clk, r781_out, r782_out);
	reg32 r783 (rst, clk, r782_out, r783_out);
	reg32 r784 (rst, clk, r783_out, r784_out);
	reg32 r785 (rst, clk, r784_out, r785_out);
	reg32 r786 (rst, clk, r785_out, r786_out);
	reg32 r787 (rst, clk, r786_out, r787_out);
	reg32 r788 (rst, clk, r787_out, r788_out);
	reg32 r789 (rst, clk, r788_out, r789_out);
	reg32 r790 (rst, clk, r789_out, r790_out);
	reg32 r791 (rst, clk, r790_out, r791_out);
	reg32 r792 (rst, clk, r791_out, r792_out);
	reg32 r793 (rst, clk, r792_out, r793_out);
	reg32 r794 (rst, clk, r793_out, r794_out);
	reg32 r795 (rst, clk, r794_out, r795_out);
	reg32 r796 (rst, clk, r795_out, r796_out);
	reg32 r797 (rst, clk, r796_out, r797_out);
	reg32 r798 (rst, clk, r797_out, r798_out);
	reg32 r799 (rst, clk, r798_out, r799_out);
	reg32 r800 (rst, clk, r799_out, r800_out);
	reg32 r801 (rst, clk, r800_out, r801_out);
	reg32 r802 (rst, clk, r801_out, r802_out);
	reg32 r803 (rst, clk, r802_out, r803_out);
	reg32 r804 (rst, clk, r803_out, r804_out);
	reg32 r805 (rst, clk, r804_out, r805_out);
	reg32 r806 (rst, clk, r805_out, r806_out);
	reg32 r807 (rst, clk, r806_out, r807_out);
	reg32 r808 (rst, clk, r807_out, r808_out);
	reg32 r809 (rst, clk, r808_out, r809_out);
	reg32 r810 (rst, clk, r809_out, r810_out);
	reg32 r811 (rst, clk, r810_out, r811_out);
	reg32 r812 (rst, clk, r811_out, r812_out);
	reg32 r813 (rst, clk, r812_out, r813_out);
	reg32 r814 (rst, clk, r813_out, r814_out);
	reg32 r815 (rst, clk, r814_out, r815_out);
	reg32 r816 (rst, clk, r815_out, r816_out);
	reg32 r817 (rst, clk, r816_out, r817_out);
	reg32 r818 (rst, clk, r817_out, r818_out);
	reg32 r819 (rst, clk, r818_out, r819_out);
	reg32 r820 (rst, clk, r819_out, r820_out);
	reg32 r821 (rst, clk, r820_out, r821_out);
	reg32 r822 (rst, clk, r821_out, r822_out);
	reg32 r823 (rst, clk, r822_out, r823_out);
	reg32 r824 (rst, clk, r823_out, r824_out);
	reg32 r825 (rst, clk, r824_out, r825_out);
	reg32 r826 (rst, clk, r825_out, r826_out);
	reg32 r827 (rst, clk, r826_out, r827_out);
	reg32 r828 (rst, clk, r827_out, r828_out);
	reg32 r829 (rst, clk, r828_out, r829_out);
	reg32 r830 (rst, clk, r829_out, r830_out);
	reg32 r831 (rst, clk, r830_out, r831_out);
	reg32 r832 (rst, clk, r831_out, r832_out);
	reg32 r833 (rst, clk, r832_out, r833_out);
	reg32 r834 (rst, clk, r833_out, r834_out);
	reg32 r835 (rst, clk, r834_out, r835_out);
	reg32 r836 (rst, clk, r835_out, r836_out);
	reg32 r837 (rst, clk, r836_out, r837_out);
	reg32 r838 (rst, clk, r837_out, r838_out);
	reg32 r839 (rst, clk, r838_out, r839_out);
	reg32 r840 (rst, clk, r839_out, r840_out);
	reg32 r841 (rst, clk, r840_out, r841_out);
	reg32 r842 (rst, clk, r841_out, r842_out);
	reg32 r843 (rst, clk, r842_out, r843_out);
	reg32 r844 (rst, clk, r843_out, r844_out);
	reg32 r845 (rst, clk, r844_out, r845_out);
	reg32 r846 (rst, clk, r845_out, r846_out);
	reg32 r847 (rst, clk, r846_out, r847_out);
	reg32 r848 (rst, clk, r847_out, r848_out);
	reg32 r849 (rst, clk, r848_out, r849_out);
	reg32 r850 (rst, clk, r849_out, r850_out);
	reg32 r851 (rst, clk, r850_out, r851_out);
	reg32 r852 (rst, clk, r851_out, r852_out);
	reg32 r853 (rst, clk, r852_out, r853_out);
	reg32 r854 (rst, clk, r853_out, r854_out);
	reg32 r855 (rst, clk, r854_out, r855_out);
	reg32 r856 (rst, clk, r855_out, r856_out);
	reg32 r857 (rst, clk, r856_out, r857_out);
	reg32 r858 (rst, clk, r857_out, r858_out);
	reg32 r859 (rst, clk, r858_out, r859_out);
	reg32 r860 (rst, clk, r859_out, r860_out);
	reg32 r861 (rst, clk, r860_out, r861_out);
	reg32 r862 (rst, clk, r861_out, r862_out);
	reg32 r863 (rst, clk, r862_out, r863_out);
	reg32 r864 (rst, clk, r863_out, r864_out);
	reg32 r865 (rst, clk, r864_out, r865_out);
	reg32 r866 (rst, clk, r865_out, r866_out);
	reg32 r867 (rst, clk, r866_out, r867_out);
	reg32 r868 (rst, clk, r867_out, r868_out);
	reg32 r869 (rst, clk, r868_out, r869_out);
	reg32 r870 (rst, clk, r869_out, r870_out);
	reg32 r871 (rst, clk, r870_out, r871_out);
	reg32 r872 (rst, clk, r871_out, r872_out);
	reg32 r873 (rst, clk, r872_out, r873_out);
	reg32 r874 (rst, clk, r873_out, r874_out);
	reg32 r875 (rst, clk, r874_out, r875_out);
	reg32 r876 (rst, clk, r875_out, r876_out);
	reg32 r877 (rst, clk, r876_out, r877_out);
	reg32 r878 (rst, clk, r877_out, r878_out);
	reg32 r879 (rst, clk, r878_out, r879_out);
	reg32 r880 (rst, clk, r879_out, r880_out);
	reg32 r881 (rst, clk, r880_out, r881_out);
	reg32 r882 (rst, clk, r881_out, r882_out);
	reg32 r883 (rst, clk, r882_out, r883_out);
	reg32 r884 (rst, clk, r883_out, r884_out);
	reg32 r885 (rst, clk, r884_out, r885_out);
	reg32 r886 (rst, clk, r885_out, r886_out);
	reg32 r887 (rst, clk, r886_out, r887_out);
	reg32 r888 (rst, clk, r887_out, r888_out);
	reg32 r889 (rst, clk, r888_out, r889_out);
	reg32 r890 (rst, clk, r889_out, r890_out);
	reg32 r891 (rst, clk, r890_out, r891_out);
	reg32 r892 (rst, clk, r891_out, r892_out);
	reg32 r893 (rst, clk, r892_out, r893_out);
	reg32 r894 (rst, clk, r893_out, r894_out);
	reg32 r895 (rst, clk, r894_out, r895_out);
	reg32 r896 (rst, clk, r895_out, r896_out);
	reg32 r897 (rst, clk, r896_out, r897_out);
	reg32 r898 (rst, clk, r897_out, r898_out);
	reg32 r899 (rst, clk, r898_out, r899_out);
	reg32 r900 (rst, clk, r899_out, r900_out);
	reg32 r901 (rst, clk, r900_out, r901_out);
	reg32 r902 (rst, clk, r901_out, r902_out);
	reg32 r903 (rst, clk, r902_out, r903_out);
	reg32 r904 (rst, clk, r903_out, r904_out);
	reg32 r905 (rst, clk, r904_out, r905_out);
	reg32 r906 (rst, clk, r905_out, r906_out);
	reg32 r907 (rst, clk, r906_out, r907_out);
	reg32 r908 (rst, clk, r907_out, r908_out);
	reg32 r909 (rst, clk, r908_out, r909_out);
	reg32 r910 (rst, clk, r909_out, r910_out);
	reg32 r911 (rst, clk, r910_out, r911_out);
	reg32 r912 (rst, clk, r911_out, r912_out);
	reg32 r913 (rst, clk, r912_out, r913_out);
	reg32 r914 (rst, clk, r913_out, r914_out);
	reg32 r915 (rst, clk, r914_out, r915_out);
	reg32 r916 (rst, clk, r915_out, r916_out);
	reg32 r917 (rst, clk, r916_out, r917_out);
	reg32 r918 (rst, clk, r917_out, r918_out);
	reg32 r919 (rst, clk, r918_out, r919_out);
	reg32 r920 (rst, clk, r919_out, r920_out);
	reg32 r921 (rst, clk, r920_out, r921_out);
	reg32 r922 (rst, clk, r921_out, r922_out);
	reg32 r923 (rst, clk, r922_out, r923_out);
	reg32 r924 (rst, clk, r923_out, r924_out);
	reg32 r925 (rst, clk, r924_out, r925_out);
	reg32 r926 (rst, clk, r925_out, r926_out);
	reg32 r927 (rst, clk, r926_out, r927_out);
	reg32 r928 (rst, clk, r927_out, r928_out);
	reg32 r929 (rst, clk, r928_out, r929_out);
	reg32 r930 (rst, clk, r929_out, r930_out);
	reg32 r931 (rst, clk, r930_out, r931_out);
	reg32 r932 (rst, clk, r931_out, r932_out);
	reg32 r933 (rst, clk, r932_out, r933_out);
	reg32 r934 (rst, clk, r933_out, r934_out);
	reg32 r935 (rst, clk, r934_out, r935_out);
	reg32 r936 (rst, clk, r935_out, r936_out);
	reg32 r937 (rst, clk, r936_out, r937_out);
	reg32 r938 (rst, clk, r937_out, r938_out);
	reg32 r939 (rst, clk, r938_out, r939_out);
	reg32 r940 (rst, clk, r939_out, r940_out);
	reg32 r941 (rst, clk, r940_out, r941_out);
	reg32 r942 (rst, clk, r941_out, r942_out);
	reg32 r943 (rst, clk, r942_out, r943_out);
	reg32 r944 (rst, clk, r943_out, r944_out);
	reg32 r945 (rst, clk, r944_out, r945_out);
	reg32 r946 (rst, clk, r945_out, r946_out);
	reg32 r947 (rst, clk, r946_out, r947_out);
	reg32 r948 (rst, clk, r947_out, r948_out);
	reg32 r949 (rst, clk, r948_out, r949_out);
	reg32 r950 (rst, clk, r949_out, r950_out);
	reg32 r951 (rst, clk, r950_out, r951_out);
	reg32 r952 (rst, clk, r951_out, r952_out);
	reg32 r953 (rst, clk, r952_out, r953_out);
	reg32 r954 (rst, clk, r953_out, r954_out);
	reg32 r955 (rst, clk, r954_out, r955_out);
	reg32 r956 (rst, clk, r955_out, r956_out);
	reg32 r957 (rst, clk, r956_out, r957_out);
	reg32 r958 (rst, clk, r957_out, r958_out);
	reg32 r959 (rst, clk, r958_out, r959_out);
	reg32 r960 (rst, clk, r959_out, r960_out);
	reg32 r961 (rst, clk, r960_out, r961_out);
	reg32 r962 (rst, clk, r961_out, r962_out);
	reg32 r963 (rst, clk, r962_out, r963_out);
	reg32 r964 (rst, clk, r963_out, r964_out);
	reg32 r965 (rst, clk, r964_out, r965_out);
	reg32 r966 (rst, clk, r965_out, r966_out);
	reg32 r967 (rst, clk, r966_out, r967_out);
	reg32 r968 (rst, clk, r967_out, r968_out);
	reg32 r969 (rst, clk, r968_out, r969_out);
	reg32 r970 (rst, clk, r969_out, r970_out);
	reg32 r971 (rst, clk, r970_out, r971_out);
	reg32 r972 (rst, clk, r971_out, r972_out);
	reg32 r973 (rst, clk, r972_out, r973_out);
	reg32 r974 (rst, clk, r973_out, r974_out);
	reg32 r975 (rst, clk, r974_out, r975_out);
	reg32 r976 (rst, clk, r975_out, r976_out);
	reg32 r977 (rst, clk, r976_out, r977_out);
	reg32 r978 (rst, clk, r977_out, r978_out);
	reg32 r979 (rst, clk, r978_out, r979_out);
	reg32 r980 (rst, clk, r979_out, r980_out);
	reg32 r981 (rst, clk, r980_out, r981_out);
	reg32 r982 (rst, clk, r981_out, r982_out);
	reg32 r983 (rst, clk, r982_out, r983_out);
	reg32 r984 (rst, clk, r983_out, r984_out);
	reg32 r985 (rst, clk, r984_out, r985_out);
	reg32 r986 (rst, clk, r985_out, r986_out);
	reg32 r987 (rst, clk, r986_out, r987_out);
	reg32 r988 (rst, clk, r987_out, r988_out);
	reg32 r989 (rst, clk, r988_out, r989_out);
	reg32 r990 (rst, clk, r989_out, r990_out);
	reg32 r991 (rst, clk, r990_out, r991_out);
	reg32 r992 (rst, clk, r991_out, r992_out);
	reg32 r993 (rst, clk, r992_out, r993_out);
	reg32 r994 (rst, clk, r993_out, r994_out);
	reg32 r995 (rst, clk, r994_out, r995_out);
	reg32 r996 (rst, clk, r995_out, r996_out);
	reg32 r997 (rst, clk, r996_out, r997_out);
	reg32 r998 (rst, clk, r997_out, r998_out);
	reg32 r999 (rst, clk, r998_out, r999_out);

	assign out = r999_out;
endmodule
