module reg3000 ( in, clk, rst, out );
	input[31:0] in;
	input clk;
	input rst;
	output[31:0] out;

	wire [31:0] r0_out;
	wire [31:0] r1_out;
	wire [31:0] r2_out;
	wire [31:0] r3_out;
	wire [31:0] r4_out;
	wire [31:0] r5_out;
	wire [31:0] r6_out;
	wire [31:0] r7_out;
	wire [31:0] r8_out;
	wire [31:0] r9_out;
	wire [31:0] r10_out;
	wire [31:0] r11_out;
	wire [31:0] r12_out;
	wire [31:0] r13_out;
	wire [31:0] r14_out;
	wire [31:0] r15_out;
	wire [31:0] r16_out;
	wire [31:0] r17_out;
	wire [31:0] r18_out;
	wire [31:0] r19_out;
	wire [31:0] r20_out;
	wire [31:0] r21_out;
	wire [31:0] r22_out;
	wire [31:0] r23_out;
	wire [31:0] r24_out;
	wire [31:0] r25_out;
	wire [31:0] r26_out;
	wire [31:0] r27_out;
	wire [31:0] r28_out;
	wire [31:0] r29_out;
	wire [31:0] r30_out;
	wire [31:0] r31_out;
	wire [31:0] r32_out;
	wire [31:0] r33_out;
	wire [31:0] r34_out;
	wire [31:0] r35_out;
	wire [31:0] r36_out;
	wire [31:0] r37_out;
	wire [31:0] r38_out;
	wire [31:0] r39_out;
	wire [31:0] r40_out;
	wire [31:0] r41_out;
	wire [31:0] r42_out;
	wire [31:0] r43_out;
	wire [31:0] r44_out;
	wire [31:0] r45_out;
	wire [31:0] r46_out;
	wire [31:0] r47_out;
	wire [31:0] r48_out;
	wire [31:0] r49_out;
	wire [31:0] r50_out;
	wire [31:0] r51_out;
	wire [31:0] r52_out;
	wire [31:0] r53_out;
	wire [31:0] r54_out;
	wire [31:0] r55_out;
	wire [31:0] r56_out;
	wire [31:0] r57_out;
	wire [31:0] r58_out;
	wire [31:0] r59_out;
	wire [31:0] r60_out;
	wire [31:0] r61_out;
	wire [31:0] r62_out;
	wire [31:0] r63_out;
	wire [31:0] r64_out;
	wire [31:0] r65_out;
	wire [31:0] r66_out;
	wire [31:0] r67_out;
	wire [31:0] r68_out;
	wire [31:0] r69_out;
	wire [31:0] r70_out;
	wire [31:0] r71_out;
	wire [31:0] r72_out;
	wire [31:0] r73_out;
	wire [31:0] r74_out;
	wire [31:0] r75_out;
	wire [31:0] r76_out;
	wire [31:0] r77_out;
	wire [31:0] r78_out;
	wire [31:0] r79_out;
	wire [31:0] r80_out;
	wire [31:0] r81_out;
	wire [31:0] r82_out;
	wire [31:0] r83_out;
	wire [31:0] r84_out;
	wire [31:0] r85_out;
	wire [31:0] r86_out;
	wire [31:0] r87_out;
	wire [31:0] r88_out;
	wire [31:0] r89_out;
	wire [31:0] r90_out;
	wire [31:0] r91_out;
	wire [31:0] r92_out;
	wire [31:0] r93_out;
	wire [31:0] r94_out;
	wire [31:0] r95_out;
	wire [31:0] r96_out;
	wire [31:0] r97_out;
	wire [31:0] r98_out;
	wire [31:0] r99_out;
	wire [31:0] r100_out;
	wire [31:0] r101_out;
	wire [31:0] r102_out;
	wire [31:0] r103_out;
	wire [31:0] r104_out;
	wire [31:0] r105_out;
	wire [31:0] r106_out;
	wire [31:0] r107_out;
	wire [31:0] r108_out;
	wire [31:0] r109_out;
	wire [31:0] r110_out;
	wire [31:0] r111_out;
	wire [31:0] r112_out;
	wire [31:0] r113_out;
	wire [31:0] r114_out;
	wire [31:0] r115_out;
	wire [31:0] r116_out;
	wire [31:0] r117_out;
	wire [31:0] r118_out;
	wire [31:0] r119_out;
	wire [31:0] r120_out;
	wire [31:0] r121_out;
	wire [31:0] r122_out;
	wire [31:0] r123_out;
	wire [31:0] r124_out;
	wire [31:0] r125_out;
	wire [31:0] r126_out;
	wire [31:0] r127_out;
	wire [31:0] r128_out;
	wire [31:0] r129_out;
	wire [31:0] r130_out;
	wire [31:0] r131_out;
	wire [31:0] r132_out;
	wire [31:0] r133_out;
	wire [31:0] r134_out;
	wire [31:0] r135_out;
	wire [31:0] r136_out;
	wire [31:0] r137_out;
	wire [31:0] r138_out;
	wire [31:0] r139_out;
	wire [31:0] r140_out;
	wire [31:0] r141_out;
	wire [31:0] r142_out;
	wire [31:0] r143_out;
	wire [31:0] r144_out;
	wire [31:0] r145_out;
	wire [31:0] r146_out;
	wire [31:0] r147_out;
	wire [31:0] r148_out;
	wire [31:0] r149_out;
	wire [31:0] r150_out;
	wire [31:0] r151_out;
	wire [31:0] r152_out;
	wire [31:0] r153_out;
	wire [31:0] r154_out;
	wire [31:0] r155_out;
	wire [31:0] r156_out;
	wire [31:0] r157_out;
	wire [31:0] r158_out;
	wire [31:0] r159_out;
	wire [31:0] r160_out;
	wire [31:0] r161_out;
	wire [31:0] r162_out;
	wire [31:0] r163_out;
	wire [31:0] r164_out;
	wire [31:0] r165_out;
	wire [31:0] r166_out;
	wire [31:0] r167_out;
	wire [31:0] r168_out;
	wire [31:0] r169_out;
	wire [31:0] r170_out;
	wire [31:0] r171_out;
	wire [31:0] r172_out;
	wire [31:0] r173_out;
	wire [31:0] r174_out;
	wire [31:0] r175_out;
	wire [31:0] r176_out;
	wire [31:0] r177_out;
	wire [31:0] r178_out;
	wire [31:0] r179_out;
	wire [31:0] r180_out;
	wire [31:0] r181_out;
	wire [31:0] r182_out;
	wire [31:0] r183_out;
	wire [31:0] r184_out;
	wire [31:0] r185_out;
	wire [31:0] r186_out;
	wire [31:0] r187_out;
	wire [31:0] r188_out;
	wire [31:0] r189_out;
	wire [31:0] r190_out;
	wire [31:0] r191_out;
	wire [31:0] r192_out;
	wire [31:0] r193_out;
	wire [31:0] r194_out;
	wire [31:0] r195_out;
	wire [31:0] r196_out;
	wire [31:0] r197_out;
	wire [31:0] r198_out;
	wire [31:0] r199_out;
	wire [31:0] r200_out;
	wire [31:0] r201_out;
	wire [31:0] r202_out;
	wire [31:0] r203_out;
	wire [31:0] r204_out;
	wire [31:0] r205_out;
	wire [31:0] r206_out;
	wire [31:0] r207_out;
	wire [31:0] r208_out;
	wire [31:0] r209_out;
	wire [31:0] r210_out;
	wire [31:0] r211_out;
	wire [31:0] r212_out;
	wire [31:0] r213_out;
	wire [31:0] r214_out;
	wire [31:0] r215_out;
	wire [31:0] r216_out;
	wire [31:0] r217_out;
	wire [31:0] r218_out;
	wire [31:0] r219_out;
	wire [31:0] r220_out;
	wire [31:0] r221_out;
	wire [31:0] r222_out;
	wire [31:0] r223_out;
	wire [31:0] r224_out;
	wire [31:0] r225_out;
	wire [31:0] r226_out;
	wire [31:0] r227_out;
	wire [31:0] r228_out;
	wire [31:0] r229_out;
	wire [31:0] r230_out;
	wire [31:0] r231_out;
	wire [31:0] r232_out;
	wire [31:0] r233_out;
	wire [31:0] r234_out;
	wire [31:0] r235_out;
	wire [31:0] r236_out;
	wire [31:0] r237_out;
	wire [31:0] r238_out;
	wire [31:0] r239_out;
	wire [31:0] r240_out;
	wire [31:0] r241_out;
	wire [31:0] r242_out;
	wire [31:0] r243_out;
	wire [31:0] r244_out;
	wire [31:0] r245_out;
	wire [31:0] r246_out;
	wire [31:0] r247_out;
	wire [31:0] r248_out;
	wire [31:0] r249_out;
	wire [31:0] r250_out;
	wire [31:0] r251_out;
	wire [31:0] r252_out;
	wire [31:0] r253_out;
	wire [31:0] r254_out;
	wire [31:0] r255_out;
	wire [31:0] r256_out;
	wire [31:0] r257_out;
	wire [31:0] r258_out;
	wire [31:0] r259_out;
	wire [31:0] r260_out;
	wire [31:0] r261_out;
	wire [31:0] r262_out;
	wire [31:0] r263_out;
	wire [31:0] r264_out;
	wire [31:0] r265_out;
	wire [31:0] r266_out;
	wire [31:0] r267_out;
	wire [31:0] r268_out;
	wire [31:0] r269_out;
	wire [31:0] r270_out;
	wire [31:0] r271_out;
	wire [31:0] r272_out;
	wire [31:0] r273_out;
	wire [31:0] r274_out;
	wire [31:0] r275_out;
	wire [31:0] r276_out;
	wire [31:0] r277_out;
	wire [31:0] r278_out;
	wire [31:0] r279_out;
	wire [31:0] r280_out;
	wire [31:0] r281_out;
	wire [31:0] r282_out;
	wire [31:0] r283_out;
	wire [31:0] r284_out;
	wire [31:0] r285_out;
	wire [31:0] r286_out;
	wire [31:0] r287_out;
	wire [31:0] r288_out;
	wire [31:0] r289_out;
	wire [31:0] r290_out;
	wire [31:0] r291_out;
	wire [31:0] r292_out;
	wire [31:0] r293_out;
	wire [31:0] r294_out;
	wire [31:0] r295_out;
	wire [31:0] r296_out;
	wire [31:0] r297_out;
	wire [31:0] r298_out;
	wire [31:0] r299_out;
	wire [31:0] r300_out;
	wire [31:0] r301_out;
	wire [31:0] r302_out;
	wire [31:0] r303_out;
	wire [31:0] r304_out;
	wire [31:0] r305_out;
	wire [31:0] r306_out;
	wire [31:0] r307_out;
	wire [31:0] r308_out;
	wire [31:0] r309_out;
	wire [31:0] r310_out;
	wire [31:0] r311_out;
	wire [31:0] r312_out;
	wire [31:0] r313_out;
	wire [31:0] r314_out;
	wire [31:0] r315_out;
	wire [31:0] r316_out;
	wire [31:0] r317_out;
	wire [31:0] r318_out;
	wire [31:0] r319_out;
	wire [31:0] r320_out;
	wire [31:0] r321_out;
	wire [31:0] r322_out;
	wire [31:0] r323_out;
	wire [31:0] r324_out;
	wire [31:0] r325_out;
	wire [31:0] r326_out;
	wire [31:0] r327_out;
	wire [31:0] r328_out;
	wire [31:0] r329_out;
	wire [31:0] r330_out;
	wire [31:0] r331_out;
	wire [31:0] r332_out;
	wire [31:0] r333_out;
	wire [31:0] r334_out;
	wire [31:0] r335_out;
	wire [31:0] r336_out;
	wire [31:0] r337_out;
	wire [31:0] r338_out;
	wire [31:0] r339_out;
	wire [31:0] r340_out;
	wire [31:0] r341_out;
	wire [31:0] r342_out;
	wire [31:0] r343_out;
	wire [31:0] r344_out;
	wire [31:0] r345_out;
	wire [31:0] r346_out;
	wire [31:0] r347_out;
	wire [31:0] r348_out;
	wire [31:0] r349_out;
	wire [31:0] r350_out;
	wire [31:0] r351_out;
	wire [31:0] r352_out;
	wire [31:0] r353_out;
	wire [31:0] r354_out;
	wire [31:0] r355_out;
	wire [31:0] r356_out;
	wire [31:0] r357_out;
	wire [31:0] r358_out;
	wire [31:0] r359_out;
	wire [31:0] r360_out;
	wire [31:0] r361_out;
	wire [31:0] r362_out;
	wire [31:0] r363_out;
	wire [31:0] r364_out;
	wire [31:0] r365_out;
	wire [31:0] r366_out;
	wire [31:0] r367_out;
	wire [31:0] r368_out;
	wire [31:0] r369_out;
	wire [31:0] r370_out;
	wire [31:0] r371_out;
	wire [31:0] r372_out;
	wire [31:0] r373_out;
	wire [31:0] r374_out;
	wire [31:0] r375_out;
	wire [31:0] r376_out;
	wire [31:0] r377_out;
	wire [31:0] r378_out;
	wire [31:0] r379_out;
	wire [31:0] r380_out;
	wire [31:0] r381_out;
	wire [31:0] r382_out;
	wire [31:0] r383_out;
	wire [31:0] r384_out;
	wire [31:0] r385_out;
	wire [31:0] r386_out;
	wire [31:0] r387_out;
	wire [31:0] r388_out;
	wire [31:0] r389_out;
	wire [31:0] r390_out;
	wire [31:0] r391_out;
	wire [31:0] r392_out;
	wire [31:0] r393_out;
	wire [31:0] r394_out;
	wire [31:0] r395_out;
	wire [31:0] r396_out;
	wire [31:0] r397_out;
	wire [31:0] r398_out;
	wire [31:0] r399_out;
	wire [31:0] r400_out;
	wire [31:0] r401_out;
	wire [31:0] r402_out;
	wire [31:0] r403_out;
	wire [31:0] r404_out;
	wire [31:0] r405_out;
	wire [31:0] r406_out;
	wire [31:0] r407_out;
	wire [31:0] r408_out;
	wire [31:0] r409_out;
	wire [31:0] r410_out;
	wire [31:0] r411_out;
	wire [31:0] r412_out;
	wire [31:0] r413_out;
	wire [31:0] r414_out;
	wire [31:0] r415_out;
	wire [31:0] r416_out;
	wire [31:0] r417_out;
	wire [31:0] r418_out;
	wire [31:0] r419_out;
	wire [31:0] r420_out;
	wire [31:0] r421_out;
	wire [31:0] r422_out;
	wire [31:0] r423_out;
	wire [31:0] r424_out;
	wire [31:0] r425_out;
	wire [31:0] r426_out;
	wire [31:0] r427_out;
	wire [31:0] r428_out;
	wire [31:0] r429_out;
	wire [31:0] r430_out;
	wire [31:0] r431_out;
	wire [31:0] r432_out;
	wire [31:0] r433_out;
	wire [31:0] r434_out;
	wire [31:0] r435_out;
	wire [31:0] r436_out;
	wire [31:0] r437_out;
	wire [31:0] r438_out;
	wire [31:0] r439_out;
	wire [31:0] r440_out;
	wire [31:0] r441_out;
	wire [31:0] r442_out;
	wire [31:0] r443_out;
	wire [31:0] r444_out;
	wire [31:0] r445_out;
	wire [31:0] r446_out;
	wire [31:0] r447_out;
	wire [31:0] r448_out;
	wire [31:0] r449_out;
	wire [31:0] r450_out;
	wire [31:0] r451_out;
	wire [31:0] r452_out;
	wire [31:0] r453_out;
	wire [31:0] r454_out;
	wire [31:0] r455_out;
	wire [31:0] r456_out;
	wire [31:0] r457_out;
	wire [31:0] r458_out;
	wire [31:0] r459_out;
	wire [31:0] r460_out;
	wire [31:0] r461_out;
	wire [31:0] r462_out;
	wire [31:0] r463_out;
	wire [31:0] r464_out;
	wire [31:0] r465_out;
	wire [31:0] r466_out;
	wire [31:0] r467_out;
	wire [31:0] r468_out;
	wire [31:0] r469_out;
	wire [31:0] r470_out;
	wire [31:0] r471_out;
	wire [31:0] r472_out;
	wire [31:0] r473_out;
	wire [31:0] r474_out;
	wire [31:0] r475_out;
	wire [31:0] r476_out;
	wire [31:0] r477_out;
	wire [31:0] r478_out;
	wire [31:0] r479_out;
	wire [31:0] r480_out;
	wire [31:0] r481_out;
	wire [31:0] r482_out;
	wire [31:0] r483_out;
	wire [31:0] r484_out;
	wire [31:0] r485_out;
	wire [31:0] r486_out;
	wire [31:0] r487_out;
	wire [31:0] r488_out;
	wire [31:0] r489_out;
	wire [31:0] r490_out;
	wire [31:0] r491_out;
	wire [31:0] r492_out;
	wire [31:0] r493_out;
	wire [31:0] r494_out;
	wire [31:0] r495_out;
	wire [31:0] r496_out;
	wire [31:0] r497_out;
	wire [31:0] r498_out;
	wire [31:0] r499_out;
	wire [31:0] r500_out;
	wire [31:0] r501_out;
	wire [31:0] r502_out;
	wire [31:0] r503_out;
	wire [31:0] r504_out;
	wire [31:0] r505_out;
	wire [31:0] r506_out;
	wire [31:0] r507_out;
	wire [31:0] r508_out;
	wire [31:0] r509_out;
	wire [31:0] r510_out;
	wire [31:0] r511_out;
	wire [31:0] r512_out;
	wire [31:0] r513_out;
	wire [31:0] r514_out;
	wire [31:0] r515_out;
	wire [31:0] r516_out;
	wire [31:0] r517_out;
	wire [31:0] r518_out;
	wire [31:0] r519_out;
	wire [31:0] r520_out;
	wire [31:0] r521_out;
	wire [31:0] r522_out;
	wire [31:0] r523_out;
	wire [31:0] r524_out;
	wire [31:0] r525_out;
	wire [31:0] r526_out;
	wire [31:0] r527_out;
	wire [31:0] r528_out;
	wire [31:0] r529_out;
	wire [31:0] r530_out;
	wire [31:0] r531_out;
	wire [31:0] r532_out;
	wire [31:0] r533_out;
	wire [31:0] r534_out;
	wire [31:0] r535_out;
	wire [31:0] r536_out;
	wire [31:0] r537_out;
	wire [31:0] r538_out;
	wire [31:0] r539_out;
	wire [31:0] r540_out;
	wire [31:0] r541_out;
	wire [31:0] r542_out;
	wire [31:0] r543_out;
	wire [31:0] r544_out;
	wire [31:0] r545_out;
	wire [31:0] r546_out;
	wire [31:0] r547_out;
	wire [31:0] r548_out;
	wire [31:0] r549_out;
	wire [31:0] r550_out;
	wire [31:0] r551_out;
	wire [31:0] r552_out;
	wire [31:0] r553_out;
	wire [31:0] r554_out;
	wire [31:0] r555_out;
	wire [31:0] r556_out;
	wire [31:0] r557_out;
	wire [31:0] r558_out;
	wire [31:0] r559_out;
	wire [31:0] r560_out;
	wire [31:0] r561_out;
	wire [31:0] r562_out;
	wire [31:0] r563_out;
	wire [31:0] r564_out;
	wire [31:0] r565_out;
	wire [31:0] r566_out;
	wire [31:0] r567_out;
	wire [31:0] r568_out;
	wire [31:0] r569_out;
	wire [31:0] r570_out;
	wire [31:0] r571_out;
	wire [31:0] r572_out;
	wire [31:0] r573_out;
	wire [31:0] r574_out;
	wire [31:0] r575_out;
	wire [31:0] r576_out;
	wire [31:0] r577_out;
	wire [31:0] r578_out;
	wire [31:0] r579_out;
	wire [31:0] r580_out;
	wire [31:0] r581_out;
	wire [31:0] r582_out;
	wire [31:0] r583_out;
	wire [31:0] r584_out;
	wire [31:0] r585_out;
	wire [31:0] r586_out;
	wire [31:0] r587_out;
	wire [31:0] r588_out;
	wire [31:0] r589_out;
	wire [31:0] r590_out;
	wire [31:0] r591_out;
	wire [31:0] r592_out;
	wire [31:0] r593_out;
	wire [31:0] r594_out;
	wire [31:0] r595_out;
	wire [31:0] r596_out;
	wire [31:0] r597_out;
	wire [31:0] r598_out;
	wire [31:0] r599_out;
	wire [31:0] r600_out;
	wire [31:0] r601_out;
	wire [31:0] r602_out;
	wire [31:0] r603_out;
	wire [31:0] r604_out;
	wire [31:0] r605_out;
	wire [31:0] r606_out;
	wire [31:0] r607_out;
	wire [31:0] r608_out;
	wire [31:0] r609_out;
	wire [31:0] r610_out;
	wire [31:0] r611_out;
	wire [31:0] r612_out;
	wire [31:0] r613_out;
	wire [31:0] r614_out;
	wire [31:0] r615_out;
	wire [31:0] r616_out;
	wire [31:0] r617_out;
	wire [31:0] r618_out;
	wire [31:0] r619_out;
	wire [31:0] r620_out;
	wire [31:0] r621_out;
	wire [31:0] r622_out;
	wire [31:0] r623_out;
	wire [31:0] r624_out;
	wire [31:0] r625_out;
	wire [31:0] r626_out;
	wire [31:0] r627_out;
	wire [31:0] r628_out;
	wire [31:0] r629_out;
	wire [31:0] r630_out;
	wire [31:0] r631_out;
	wire [31:0] r632_out;
	wire [31:0] r633_out;
	wire [31:0] r634_out;
	wire [31:0] r635_out;
	wire [31:0] r636_out;
	wire [31:0] r637_out;
	wire [31:0] r638_out;
	wire [31:0] r639_out;
	wire [31:0] r640_out;
	wire [31:0] r641_out;
	wire [31:0] r642_out;
	wire [31:0] r643_out;
	wire [31:0] r644_out;
	wire [31:0] r645_out;
	wire [31:0] r646_out;
	wire [31:0] r647_out;
	wire [31:0] r648_out;
	wire [31:0] r649_out;
	wire [31:0] r650_out;
	wire [31:0] r651_out;
	wire [31:0] r652_out;
	wire [31:0] r653_out;
	wire [31:0] r654_out;
	wire [31:0] r655_out;
	wire [31:0] r656_out;
	wire [31:0] r657_out;
	wire [31:0] r658_out;
	wire [31:0] r659_out;
	wire [31:0] r660_out;
	wire [31:0] r661_out;
	wire [31:0] r662_out;
	wire [31:0] r663_out;
	wire [31:0] r664_out;
	wire [31:0] r665_out;
	wire [31:0] r666_out;
	wire [31:0] r667_out;
	wire [31:0] r668_out;
	wire [31:0] r669_out;
	wire [31:0] r670_out;
	wire [31:0] r671_out;
	wire [31:0] r672_out;
	wire [31:0] r673_out;
	wire [31:0] r674_out;
	wire [31:0] r675_out;
	wire [31:0] r676_out;
	wire [31:0] r677_out;
	wire [31:0] r678_out;
	wire [31:0] r679_out;
	wire [31:0] r680_out;
	wire [31:0] r681_out;
	wire [31:0] r682_out;
	wire [31:0] r683_out;
	wire [31:0] r684_out;
	wire [31:0] r685_out;
	wire [31:0] r686_out;
	wire [31:0] r687_out;
	wire [31:0] r688_out;
	wire [31:0] r689_out;
	wire [31:0] r690_out;
	wire [31:0] r691_out;
	wire [31:0] r692_out;
	wire [31:0] r693_out;
	wire [31:0] r694_out;
	wire [31:0] r695_out;
	wire [31:0] r696_out;
	wire [31:0] r697_out;
	wire [31:0] r698_out;
	wire [31:0] r699_out;
	wire [31:0] r700_out;
	wire [31:0] r701_out;
	wire [31:0] r702_out;
	wire [31:0] r703_out;
	wire [31:0] r704_out;
	wire [31:0] r705_out;
	wire [31:0] r706_out;
	wire [31:0] r707_out;
	wire [31:0] r708_out;
	wire [31:0] r709_out;
	wire [31:0] r710_out;
	wire [31:0] r711_out;
	wire [31:0] r712_out;
	wire [31:0] r713_out;
	wire [31:0] r714_out;
	wire [31:0] r715_out;
	wire [31:0] r716_out;
	wire [31:0] r717_out;
	wire [31:0] r718_out;
	wire [31:0] r719_out;
	wire [31:0] r720_out;
	wire [31:0] r721_out;
	wire [31:0] r722_out;
	wire [31:0] r723_out;
	wire [31:0] r724_out;
	wire [31:0] r725_out;
	wire [31:0] r726_out;
	wire [31:0] r727_out;
	wire [31:0] r728_out;
	wire [31:0] r729_out;
	wire [31:0] r730_out;
	wire [31:0] r731_out;
	wire [31:0] r732_out;
	wire [31:0] r733_out;
	wire [31:0] r734_out;
	wire [31:0] r735_out;
	wire [31:0] r736_out;
	wire [31:0] r737_out;
	wire [31:0] r738_out;
	wire [31:0] r739_out;
	wire [31:0] r740_out;
	wire [31:0] r741_out;
	wire [31:0] r742_out;
	wire [31:0] r743_out;
	wire [31:0] r744_out;
	wire [31:0] r745_out;
	wire [31:0] r746_out;
	wire [31:0] r747_out;
	wire [31:0] r748_out;
	wire [31:0] r749_out;
	wire [31:0] r750_out;
	wire [31:0] r751_out;
	wire [31:0] r752_out;
	wire [31:0] r753_out;
	wire [31:0] r754_out;
	wire [31:0] r755_out;
	wire [31:0] r756_out;
	wire [31:0] r757_out;
	wire [31:0] r758_out;
	wire [31:0] r759_out;
	wire [31:0] r760_out;
	wire [31:0] r761_out;
	wire [31:0] r762_out;
	wire [31:0] r763_out;
	wire [31:0] r764_out;
	wire [31:0] r765_out;
	wire [31:0] r766_out;
	wire [31:0] r767_out;
	wire [31:0] r768_out;
	wire [31:0] r769_out;
	wire [31:0] r770_out;
	wire [31:0] r771_out;
	wire [31:0] r772_out;
	wire [31:0] r773_out;
	wire [31:0] r774_out;
	wire [31:0] r775_out;
	wire [31:0] r776_out;
	wire [31:0] r777_out;
	wire [31:0] r778_out;
	wire [31:0] r779_out;
	wire [31:0] r780_out;
	wire [31:0] r781_out;
	wire [31:0] r782_out;
	wire [31:0] r783_out;
	wire [31:0] r784_out;
	wire [31:0] r785_out;
	wire [31:0] r786_out;
	wire [31:0] r787_out;
	wire [31:0] r788_out;
	wire [31:0] r789_out;
	wire [31:0] r790_out;
	wire [31:0] r791_out;
	wire [31:0] r792_out;
	wire [31:0] r793_out;
	wire [31:0] r794_out;
	wire [31:0] r795_out;
	wire [31:0] r796_out;
	wire [31:0] r797_out;
	wire [31:0] r798_out;
	wire [31:0] r799_out;
	wire [31:0] r800_out;
	wire [31:0] r801_out;
	wire [31:0] r802_out;
	wire [31:0] r803_out;
	wire [31:0] r804_out;
	wire [31:0] r805_out;
	wire [31:0] r806_out;
	wire [31:0] r807_out;
	wire [31:0] r808_out;
	wire [31:0] r809_out;
	wire [31:0] r810_out;
	wire [31:0] r811_out;
	wire [31:0] r812_out;
	wire [31:0] r813_out;
	wire [31:0] r814_out;
	wire [31:0] r815_out;
	wire [31:0] r816_out;
	wire [31:0] r817_out;
	wire [31:0] r818_out;
	wire [31:0] r819_out;
	wire [31:0] r820_out;
	wire [31:0] r821_out;
	wire [31:0] r822_out;
	wire [31:0] r823_out;
	wire [31:0] r824_out;
	wire [31:0] r825_out;
	wire [31:0] r826_out;
	wire [31:0] r827_out;
	wire [31:0] r828_out;
	wire [31:0] r829_out;
	wire [31:0] r830_out;
	wire [31:0] r831_out;
	wire [31:0] r832_out;
	wire [31:0] r833_out;
	wire [31:0] r834_out;
	wire [31:0] r835_out;
	wire [31:0] r836_out;
	wire [31:0] r837_out;
	wire [31:0] r838_out;
	wire [31:0] r839_out;
	wire [31:0] r840_out;
	wire [31:0] r841_out;
	wire [31:0] r842_out;
	wire [31:0] r843_out;
	wire [31:0] r844_out;
	wire [31:0] r845_out;
	wire [31:0] r846_out;
	wire [31:0] r847_out;
	wire [31:0] r848_out;
	wire [31:0] r849_out;
	wire [31:0] r850_out;
	wire [31:0] r851_out;
	wire [31:0] r852_out;
	wire [31:0] r853_out;
	wire [31:0] r854_out;
	wire [31:0] r855_out;
	wire [31:0] r856_out;
	wire [31:0] r857_out;
	wire [31:0] r858_out;
	wire [31:0] r859_out;
	wire [31:0] r860_out;
	wire [31:0] r861_out;
	wire [31:0] r862_out;
	wire [31:0] r863_out;
	wire [31:0] r864_out;
	wire [31:0] r865_out;
	wire [31:0] r866_out;
	wire [31:0] r867_out;
	wire [31:0] r868_out;
	wire [31:0] r869_out;
	wire [31:0] r870_out;
	wire [31:0] r871_out;
	wire [31:0] r872_out;
	wire [31:0] r873_out;
	wire [31:0] r874_out;
	wire [31:0] r875_out;
	wire [31:0] r876_out;
	wire [31:0] r877_out;
	wire [31:0] r878_out;
	wire [31:0] r879_out;
	wire [31:0] r880_out;
	wire [31:0] r881_out;
	wire [31:0] r882_out;
	wire [31:0] r883_out;
	wire [31:0] r884_out;
	wire [31:0] r885_out;
	wire [31:0] r886_out;
	wire [31:0] r887_out;
	wire [31:0] r888_out;
	wire [31:0] r889_out;
	wire [31:0] r890_out;
	wire [31:0] r891_out;
	wire [31:0] r892_out;
	wire [31:0] r893_out;
	wire [31:0] r894_out;
	wire [31:0] r895_out;
	wire [31:0] r896_out;
	wire [31:0] r897_out;
	wire [31:0] r898_out;
	wire [31:0] r899_out;
	wire [31:0] r900_out;
	wire [31:0] r901_out;
	wire [31:0] r902_out;
	wire [31:0] r903_out;
	wire [31:0] r904_out;
	wire [31:0] r905_out;
	wire [31:0] r906_out;
	wire [31:0] r907_out;
	wire [31:0] r908_out;
	wire [31:0] r909_out;
	wire [31:0] r910_out;
	wire [31:0] r911_out;
	wire [31:0] r912_out;
	wire [31:0] r913_out;
	wire [31:0] r914_out;
	wire [31:0] r915_out;
	wire [31:0] r916_out;
	wire [31:0] r917_out;
	wire [31:0] r918_out;
	wire [31:0] r919_out;
	wire [31:0] r920_out;
	wire [31:0] r921_out;
	wire [31:0] r922_out;
	wire [31:0] r923_out;
	wire [31:0] r924_out;
	wire [31:0] r925_out;
	wire [31:0] r926_out;
	wire [31:0] r927_out;
	wire [31:0] r928_out;
	wire [31:0] r929_out;
	wire [31:0] r930_out;
	wire [31:0] r931_out;
	wire [31:0] r932_out;
	wire [31:0] r933_out;
	wire [31:0] r934_out;
	wire [31:0] r935_out;
	wire [31:0] r936_out;
	wire [31:0] r937_out;
	wire [31:0] r938_out;
	wire [31:0] r939_out;
	wire [31:0] r940_out;
	wire [31:0] r941_out;
	wire [31:0] r942_out;
	wire [31:0] r943_out;
	wire [31:0] r944_out;
	wire [31:0] r945_out;
	wire [31:0] r946_out;
	wire [31:0] r947_out;
	wire [31:0] r948_out;
	wire [31:0] r949_out;
	wire [31:0] r950_out;
	wire [31:0] r951_out;
	wire [31:0] r952_out;
	wire [31:0] r953_out;
	wire [31:0] r954_out;
	wire [31:0] r955_out;
	wire [31:0] r956_out;
	wire [31:0] r957_out;
	wire [31:0] r958_out;
	wire [31:0] r959_out;
	wire [31:0] r960_out;
	wire [31:0] r961_out;
	wire [31:0] r962_out;
	wire [31:0] r963_out;
	wire [31:0] r964_out;
	wire [31:0] r965_out;
	wire [31:0] r966_out;
	wire [31:0] r967_out;
	wire [31:0] r968_out;
	wire [31:0] r969_out;
	wire [31:0] r970_out;
	wire [31:0] r971_out;
	wire [31:0] r972_out;
	wire [31:0] r973_out;
	wire [31:0] r974_out;
	wire [31:0] r975_out;
	wire [31:0] r976_out;
	wire [31:0] r977_out;
	wire [31:0] r978_out;
	wire [31:0] r979_out;
	wire [31:0] r980_out;
	wire [31:0] r981_out;
	wire [31:0] r982_out;
	wire [31:0] r983_out;
	wire [31:0] r984_out;
	wire [31:0] r985_out;
	wire [31:0] r986_out;
	wire [31:0] r987_out;
	wire [31:0] r988_out;
	wire [31:0] r989_out;
	wire [31:0] r990_out;
	wire [31:0] r991_out;
	wire [31:0] r992_out;
	wire [31:0] r993_out;
	wire [31:0] r994_out;
	wire [31:0] r995_out;
	wire [31:0] r996_out;
	wire [31:0] r997_out;
	wire [31:0] r998_out;
	wire [31:0] r999_out;
	wire [31:0] r1000_out;
	wire [31:0] r1001_out;
	wire [31:0] r1002_out;
	wire [31:0] r1003_out;
	wire [31:0] r1004_out;
	wire [31:0] r1005_out;
	wire [31:0] r1006_out;
	wire [31:0] r1007_out;
	wire [31:0] r1008_out;
	wire [31:0] r1009_out;
	wire [31:0] r1010_out;
	wire [31:0] r1011_out;
	wire [31:0] r1012_out;
	wire [31:0] r1013_out;
	wire [31:0] r1014_out;
	wire [31:0] r1015_out;
	wire [31:0] r1016_out;
	wire [31:0] r1017_out;
	wire [31:0] r1018_out;
	wire [31:0] r1019_out;
	wire [31:0] r1020_out;
	wire [31:0] r1021_out;
	wire [31:0] r1022_out;
	wire [31:0] r1023_out;
	wire [31:0] r1024_out;
	wire [31:0] r1025_out;
	wire [31:0] r1026_out;
	wire [31:0] r1027_out;
	wire [31:0] r1028_out;
	wire [31:0] r1029_out;
	wire [31:0] r1030_out;
	wire [31:0] r1031_out;
	wire [31:0] r1032_out;
	wire [31:0] r1033_out;
	wire [31:0] r1034_out;
	wire [31:0] r1035_out;
	wire [31:0] r1036_out;
	wire [31:0] r1037_out;
	wire [31:0] r1038_out;
	wire [31:0] r1039_out;
	wire [31:0] r1040_out;
	wire [31:0] r1041_out;
	wire [31:0] r1042_out;
	wire [31:0] r1043_out;
	wire [31:0] r1044_out;
	wire [31:0] r1045_out;
	wire [31:0] r1046_out;
	wire [31:0] r1047_out;
	wire [31:0] r1048_out;
	wire [31:0] r1049_out;
	wire [31:0] r1050_out;
	wire [31:0] r1051_out;
	wire [31:0] r1052_out;
	wire [31:0] r1053_out;
	wire [31:0] r1054_out;
	wire [31:0] r1055_out;
	wire [31:0] r1056_out;
	wire [31:0] r1057_out;
	wire [31:0] r1058_out;
	wire [31:0] r1059_out;
	wire [31:0] r1060_out;
	wire [31:0] r1061_out;
	wire [31:0] r1062_out;
	wire [31:0] r1063_out;
	wire [31:0] r1064_out;
	wire [31:0] r1065_out;
	wire [31:0] r1066_out;
	wire [31:0] r1067_out;
	wire [31:0] r1068_out;
	wire [31:0] r1069_out;
	wire [31:0] r1070_out;
	wire [31:0] r1071_out;
	wire [31:0] r1072_out;
	wire [31:0] r1073_out;
	wire [31:0] r1074_out;
	wire [31:0] r1075_out;
	wire [31:0] r1076_out;
	wire [31:0] r1077_out;
	wire [31:0] r1078_out;
	wire [31:0] r1079_out;
	wire [31:0] r1080_out;
	wire [31:0] r1081_out;
	wire [31:0] r1082_out;
	wire [31:0] r1083_out;
	wire [31:0] r1084_out;
	wire [31:0] r1085_out;
	wire [31:0] r1086_out;
	wire [31:0] r1087_out;
	wire [31:0] r1088_out;
	wire [31:0] r1089_out;
	wire [31:0] r1090_out;
	wire [31:0] r1091_out;
	wire [31:0] r1092_out;
	wire [31:0] r1093_out;
	wire [31:0] r1094_out;
	wire [31:0] r1095_out;
	wire [31:0] r1096_out;
	wire [31:0] r1097_out;
	wire [31:0] r1098_out;
	wire [31:0] r1099_out;
	wire [31:0] r1100_out;
	wire [31:0] r1101_out;
	wire [31:0] r1102_out;
	wire [31:0] r1103_out;
	wire [31:0] r1104_out;
	wire [31:0] r1105_out;
	wire [31:0] r1106_out;
	wire [31:0] r1107_out;
	wire [31:0] r1108_out;
	wire [31:0] r1109_out;
	wire [31:0] r1110_out;
	wire [31:0] r1111_out;
	wire [31:0] r1112_out;
	wire [31:0] r1113_out;
	wire [31:0] r1114_out;
	wire [31:0] r1115_out;
	wire [31:0] r1116_out;
	wire [31:0] r1117_out;
	wire [31:0] r1118_out;
	wire [31:0] r1119_out;
	wire [31:0] r1120_out;
	wire [31:0] r1121_out;
	wire [31:0] r1122_out;
	wire [31:0] r1123_out;
	wire [31:0] r1124_out;
	wire [31:0] r1125_out;
	wire [31:0] r1126_out;
	wire [31:0] r1127_out;
	wire [31:0] r1128_out;
	wire [31:0] r1129_out;
	wire [31:0] r1130_out;
	wire [31:0] r1131_out;
	wire [31:0] r1132_out;
	wire [31:0] r1133_out;
	wire [31:0] r1134_out;
	wire [31:0] r1135_out;
	wire [31:0] r1136_out;
	wire [31:0] r1137_out;
	wire [31:0] r1138_out;
	wire [31:0] r1139_out;
	wire [31:0] r1140_out;
	wire [31:0] r1141_out;
	wire [31:0] r1142_out;
	wire [31:0] r1143_out;
	wire [31:0] r1144_out;
	wire [31:0] r1145_out;
	wire [31:0] r1146_out;
	wire [31:0] r1147_out;
	wire [31:0] r1148_out;
	wire [31:0] r1149_out;
	wire [31:0] r1150_out;
	wire [31:0] r1151_out;
	wire [31:0] r1152_out;
	wire [31:0] r1153_out;
	wire [31:0] r1154_out;
	wire [31:0] r1155_out;
	wire [31:0] r1156_out;
	wire [31:0] r1157_out;
	wire [31:0] r1158_out;
	wire [31:0] r1159_out;
	wire [31:0] r1160_out;
	wire [31:0] r1161_out;
	wire [31:0] r1162_out;
	wire [31:0] r1163_out;
	wire [31:0] r1164_out;
	wire [31:0] r1165_out;
	wire [31:0] r1166_out;
	wire [31:0] r1167_out;
	wire [31:0] r1168_out;
	wire [31:0] r1169_out;
	wire [31:0] r1170_out;
	wire [31:0] r1171_out;
	wire [31:0] r1172_out;
	wire [31:0] r1173_out;
	wire [31:0] r1174_out;
	wire [31:0] r1175_out;
	wire [31:0] r1176_out;
	wire [31:0] r1177_out;
	wire [31:0] r1178_out;
	wire [31:0] r1179_out;
	wire [31:0] r1180_out;
	wire [31:0] r1181_out;
	wire [31:0] r1182_out;
	wire [31:0] r1183_out;
	wire [31:0] r1184_out;
	wire [31:0] r1185_out;
	wire [31:0] r1186_out;
	wire [31:0] r1187_out;
	wire [31:0] r1188_out;
	wire [31:0] r1189_out;
	wire [31:0] r1190_out;
	wire [31:0] r1191_out;
	wire [31:0] r1192_out;
	wire [31:0] r1193_out;
	wire [31:0] r1194_out;
	wire [31:0] r1195_out;
	wire [31:0] r1196_out;
	wire [31:0] r1197_out;
	wire [31:0] r1198_out;
	wire [31:0] r1199_out;
	wire [31:0] r1200_out;
	wire [31:0] r1201_out;
	wire [31:0] r1202_out;
	wire [31:0] r1203_out;
	wire [31:0] r1204_out;
	wire [31:0] r1205_out;
	wire [31:0] r1206_out;
	wire [31:0] r1207_out;
	wire [31:0] r1208_out;
	wire [31:0] r1209_out;
	wire [31:0] r1210_out;
	wire [31:0] r1211_out;
	wire [31:0] r1212_out;
	wire [31:0] r1213_out;
	wire [31:0] r1214_out;
	wire [31:0] r1215_out;
	wire [31:0] r1216_out;
	wire [31:0] r1217_out;
	wire [31:0] r1218_out;
	wire [31:0] r1219_out;
	wire [31:0] r1220_out;
	wire [31:0] r1221_out;
	wire [31:0] r1222_out;
	wire [31:0] r1223_out;
	wire [31:0] r1224_out;
	wire [31:0] r1225_out;
	wire [31:0] r1226_out;
	wire [31:0] r1227_out;
	wire [31:0] r1228_out;
	wire [31:0] r1229_out;
	wire [31:0] r1230_out;
	wire [31:0] r1231_out;
	wire [31:0] r1232_out;
	wire [31:0] r1233_out;
	wire [31:0] r1234_out;
	wire [31:0] r1235_out;
	wire [31:0] r1236_out;
	wire [31:0] r1237_out;
	wire [31:0] r1238_out;
	wire [31:0] r1239_out;
	wire [31:0] r1240_out;
	wire [31:0] r1241_out;
	wire [31:0] r1242_out;
	wire [31:0] r1243_out;
	wire [31:0] r1244_out;
	wire [31:0] r1245_out;
	wire [31:0] r1246_out;
	wire [31:0] r1247_out;
	wire [31:0] r1248_out;
	wire [31:0] r1249_out;
	wire [31:0] r1250_out;
	wire [31:0] r1251_out;
	wire [31:0] r1252_out;
	wire [31:0] r1253_out;
	wire [31:0] r1254_out;
	wire [31:0] r1255_out;
	wire [31:0] r1256_out;
	wire [31:0] r1257_out;
	wire [31:0] r1258_out;
	wire [31:0] r1259_out;
	wire [31:0] r1260_out;
	wire [31:0] r1261_out;
	wire [31:0] r1262_out;
	wire [31:0] r1263_out;
	wire [31:0] r1264_out;
	wire [31:0] r1265_out;
	wire [31:0] r1266_out;
	wire [31:0] r1267_out;
	wire [31:0] r1268_out;
	wire [31:0] r1269_out;
	wire [31:0] r1270_out;
	wire [31:0] r1271_out;
	wire [31:0] r1272_out;
	wire [31:0] r1273_out;
	wire [31:0] r1274_out;
	wire [31:0] r1275_out;
	wire [31:0] r1276_out;
	wire [31:0] r1277_out;
	wire [31:0] r1278_out;
	wire [31:0] r1279_out;
	wire [31:0] r1280_out;
	wire [31:0] r1281_out;
	wire [31:0] r1282_out;
	wire [31:0] r1283_out;
	wire [31:0] r1284_out;
	wire [31:0] r1285_out;
	wire [31:0] r1286_out;
	wire [31:0] r1287_out;
	wire [31:0] r1288_out;
	wire [31:0] r1289_out;
	wire [31:0] r1290_out;
	wire [31:0] r1291_out;
	wire [31:0] r1292_out;
	wire [31:0] r1293_out;
	wire [31:0] r1294_out;
	wire [31:0] r1295_out;
	wire [31:0] r1296_out;
	wire [31:0] r1297_out;
	wire [31:0] r1298_out;
	wire [31:0] r1299_out;
	wire [31:0] r1300_out;
	wire [31:0] r1301_out;
	wire [31:0] r1302_out;
	wire [31:0] r1303_out;
	wire [31:0] r1304_out;
	wire [31:0] r1305_out;
	wire [31:0] r1306_out;
	wire [31:0] r1307_out;
	wire [31:0] r1308_out;
	wire [31:0] r1309_out;
	wire [31:0] r1310_out;
	wire [31:0] r1311_out;
	wire [31:0] r1312_out;
	wire [31:0] r1313_out;
	wire [31:0] r1314_out;
	wire [31:0] r1315_out;
	wire [31:0] r1316_out;
	wire [31:0] r1317_out;
	wire [31:0] r1318_out;
	wire [31:0] r1319_out;
	wire [31:0] r1320_out;
	wire [31:0] r1321_out;
	wire [31:0] r1322_out;
	wire [31:0] r1323_out;
	wire [31:0] r1324_out;
	wire [31:0] r1325_out;
	wire [31:0] r1326_out;
	wire [31:0] r1327_out;
	wire [31:0] r1328_out;
	wire [31:0] r1329_out;
	wire [31:0] r1330_out;
	wire [31:0] r1331_out;
	wire [31:0] r1332_out;
	wire [31:0] r1333_out;
	wire [31:0] r1334_out;
	wire [31:0] r1335_out;
	wire [31:0] r1336_out;
	wire [31:0] r1337_out;
	wire [31:0] r1338_out;
	wire [31:0] r1339_out;
	wire [31:0] r1340_out;
	wire [31:0] r1341_out;
	wire [31:0] r1342_out;
	wire [31:0] r1343_out;
	wire [31:0] r1344_out;
	wire [31:0] r1345_out;
	wire [31:0] r1346_out;
	wire [31:0] r1347_out;
	wire [31:0] r1348_out;
	wire [31:0] r1349_out;
	wire [31:0] r1350_out;
	wire [31:0] r1351_out;
	wire [31:0] r1352_out;
	wire [31:0] r1353_out;
	wire [31:0] r1354_out;
	wire [31:0] r1355_out;
	wire [31:0] r1356_out;
	wire [31:0] r1357_out;
	wire [31:0] r1358_out;
	wire [31:0] r1359_out;
	wire [31:0] r1360_out;
	wire [31:0] r1361_out;
	wire [31:0] r1362_out;
	wire [31:0] r1363_out;
	wire [31:0] r1364_out;
	wire [31:0] r1365_out;
	wire [31:0] r1366_out;
	wire [31:0] r1367_out;
	wire [31:0] r1368_out;
	wire [31:0] r1369_out;
	wire [31:0] r1370_out;
	wire [31:0] r1371_out;
	wire [31:0] r1372_out;
	wire [31:0] r1373_out;
	wire [31:0] r1374_out;
	wire [31:0] r1375_out;
	wire [31:0] r1376_out;
	wire [31:0] r1377_out;
	wire [31:0] r1378_out;
	wire [31:0] r1379_out;
	wire [31:0] r1380_out;
	wire [31:0] r1381_out;
	wire [31:0] r1382_out;
	wire [31:0] r1383_out;
	wire [31:0] r1384_out;
	wire [31:0] r1385_out;
	wire [31:0] r1386_out;
	wire [31:0] r1387_out;
	wire [31:0] r1388_out;
	wire [31:0] r1389_out;
	wire [31:0] r1390_out;
	wire [31:0] r1391_out;
	wire [31:0] r1392_out;
	wire [31:0] r1393_out;
	wire [31:0] r1394_out;
	wire [31:0] r1395_out;
	wire [31:0] r1396_out;
	wire [31:0] r1397_out;
	wire [31:0] r1398_out;
	wire [31:0] r1399_out;
	wire [31:0] r1400_out;
	wire [31:0] r1401_out;
	wire [31:0] r1402_out;
	wire [31:0] r1403_out;
	wire [31:0] r1404_out;
	wire [31:0] r1405_out;
	wire [31:0] r1406_out;
	wire [31:0] r1407_out;
	wire [31:0] r1408_out;
	wire [31:0] r1409_out;
	wire [31:0] r1410_out;
	wire [31:0] r1411_out;
	wire [31:0] r1412_out;
	wire [31:0] r1413_out;
	wire [31:0] r1414_out;
	wire [31:0] r1415_out;
	wire [31:0] r1416_out;
	wire [31:0] r1417_out;
	wire [31:0] r1418_out;
	wire [31:0] r1419_out;
	wire [31:0] r1420_out;
	wire [31:0] r1421_out;
	wire [31:0] r1422_out;
	wire [31:0] r1423_out;
	wire [31:0] r1424_out;
	wire [31:0] r1425_out;
	wire [31:0] r1426_out;
	wire [31:0] r1427_out;
	wire [31:0] r1428_out;
	wire [31:0] r1429_out;
	wire [31:0] r1430_out;
	wire [31:0] r1431_out;
	wire [31:0] r1432_out;
	wire [31:0] r1433_out;
	wire [31:0] r1434_out;
	wire [31:0] r1435_out;
	wire [31:0] r1436_out;
	wire [31:0] r1437_out;
	wire [31:0] r1438_out;
	wire [31:0] r1439_out;
	wire [31:0] r1440_out;
	wire [31:0] r1441_out;
	wire [31:0] r1442_out;
	wire [31:0] r1443_out;
	wire [31:0] r1444_out;
	wire [31:0] r1445_out;
	wire [31:0] r1446_out;
	wire [31:0] r1447_out;
	wire [31:0] r1448_out;
	wire [31:0] r1449_out;
	wire [31:0] r1450_out;
	wire [31:0] r1451_out;
	wire [31:0] r1452_out;
	wire [31:0] r1453_out;
	wire [31:0] r1454_out;
	wire [31:0] r1455_out;
	wire [31:0] r1456_out;
	wire [31:0] r1457_out;
	wire [31:0] r1458_out;
	wire [31:0] r1459_out;
	wire [31:0] r1460_out;
	wire [31:0] r1461_out;
	wire [31:0] r1462_out;
	wire [31:0] r1463_out;
	wire [31:0] r1464_out;
	wire [31:0] r1465_out;
	wire [31:0] r1466_out;
	wire [31:0] r1467_out;
	wire [31:0] r1468_out;
	wire [31:0] r1469_out;
	wire [31:0] r1470_out;
	wire [31:0] r1471_out;
	wire [31:0] r1472_out;
	wire [31:0] r1473_out;
	wire [31:0] r1474_out;
	wire [31:0] r1475_out;
	wire [31:0] r1476_out;
	wire [31:0] r1477_out;
	wire [31:0] r1478_out;
	wire [31:0] r1479_out;
	wire [31:0] r1480_out;
	wire [31:0] r1481_out;
	wire [31:0] r1482_out;
	wire [31:0] r1483_out;
	wire [31:0] r1484_out;
	wire [31:0] r1485_out;
	wire [31:0] r1486_out;
	wire [31:0] r1487_out;
	wire [31:0] r1488_out;
	wire [31:0] r1489_out;
	wire [31:0] r1490_out;
	wire [31:0] r1491_out;
	wire [31:0] r1492_out;
	wire [31:0] r1493_out;
	wire [31:0] r1494_out;
	wire [31:0] r1495_out;
	wire [31:0] r1496_out;
	wire [31:0] r1497_out;
	wire [31:0] r1498_out;
	wire [31:0] r1499_out;
	wire [31:0] r1500_out;
	wire [31:0] r1501_out;
	wire [31:0] r1502_out;
	wire [31:0] r1503_out;
	wire [31:0] r1504_out;
	wire [31:0] r1505_out;
	wire [31:0] r1506_out;
	wire [31:0] r1507_out;
	wire [31:0] r1508_out;
	wire [31:0] r1509_out;
	wire [31:0] r1510_out;
	wire [31:0] r1511_out;
	wire [31:0] r1512_out;
	wire [31:0] r1513_out;
	wire [31:0] r1514_out;
	wire [31:0] r1515_out;
	wire [31:0] r1516_out;
	wire [31:0] r1517_out;
	wire [31:0] r1518_out;
	wire [31:0] r1519_out;
	wire [31:0] r1520_out;
	wire [31:0] r1521_out;
	wire [31:0] r1522_out;
	wire [31:0] r1523_out;
	wire [31:0] r1524_out;
	wire [31:0] r1525_out;
	wire [31:0] r1526_out;
	wire [31:0] r1527_out;
	wire [31:0] r1528_out;
	wire [31:0] r1529_out;
	wire [31:0] r1530_out;
	wire [31:0] r1531_out;
	wire [31:0] r1532_out;
	wire [31:0] r1533_out;
	wire [31:0] r1534_out;
	wire [31:0] r1535_out;
	wire [31:0] r1536_out;
	wire [31:0] r1537_out;
	wire [31:0] r1538_out;
	wire [31:0] r1539_out;
	wire [31:0] r1540_out;
	wire [31:0] r1541_out;
	wire [31:0] r1542_out;
	wire [31:0] r1543_out;
	wire [31:0] r1544_out;
	wire [31:0] r1545_out;
	wire [31:0] r1546_out;
	wire [31:0] r1547_out;
	wire [31:0] r1548_out;
	wire [31:0] r1549_out;
	wire [31:0] r1550_out;
	wire [31:0] r1551_out;
	wire [31:0] r1552_out;
	wire [31:0] r1553_out;
	wire [31:0] r1554_out;
	wire [31:0] r1555_out;
	wire [31:0] r1556_out;
	wire [31:0] r1557_out;
	wire [31:0] r1558_out;
	wire [31:0] r1559_out;
	wire [31:0] r1560_out;
	wire [31:0] r1561_out;
	wire [31:0] r1562_out;
	wire [31:0] r1563_out;
	wire [31:0] r1564_out;
	wire [31:0] r1565_out;
	wire [31:0] r1566_out;
	wire [31:0] r1567_out;
	wire [31:0] r1568_out;
	wire [31:0] r1569_out;
	wire [31:0] r1570_out;
	wire [31:0] r1571_out;
	wire [31:0] r1572_out;
	wire [31:0] r1573_out;
	wire [31:0] r1574_out;
	wire [31:0] r1575_out;
	wire [31:0] r1576_out;
	wire [31:0] r1577_out;
	wire [31:0] r1578_out;
	wire [31:0] r1579_out;
	wire [31:0] r1580_out;
	wire [31:0] r1581_out;
	wire [31:0] r1582_out;
	wire [31:0] r1583_out;
	wire [31:0] r1584_out;
	wire [31:0] r1585_out;
	wire [31:0] r1586_out;
	wire [31:0] r1587_out;
	wire [31:0] r1588_out;
	wire [31:0] r1589_out;
	wire [31:0] r1590_out;
	wire [31:0] r1591_out;
	wire [31:0] r1592_out;
	wire [31:0] r1593_out;
	wire [31:0] r1594_out;
	wire [31:0] r1595_out;
	wire [31:0] r1596_out;
	wire [31:0] r1597_out;
	wire [31:0] r1598_out;
	wire [31:0] r1599_out;
	wire [31:0] r1600_out;
	wire [31:0] r1601_out;
	wire [31:0] r1602_out;
	wire [31:0] r1603_out;
	wire [31:0] r1604_out;
	wire [31:0] r1605_out;
	wire [31:0] r1606_out;
	wire [31:0] r1607_out;
	wire [31:0] r1608_out;
	wire [31:0] r1609_out;
	wire [31:0] r1610_out;
	wire [31:0] r1611_out;
	wire [31:0] r1612_out;
	wire [31:0] r1613_out;
	wire [31:0] r1614_out;
	wire [31:0] r1615_out;
	wire [31:0] r1616_out;
	wire [31:0] r1617_out;
	wire [31:0] r1618_out;
	wire [31:0] r1619_out;
	wire [31:0] r1620_out;
	wire [31:0] r1621_out;
	wire [31:0] r1622_out;
	wire [31:0] r1623_out;
	wire [31:0] r1624_out;
	wire [31:0] r1625_out;
	wire [31:0] r1626_out;
	wire [31:0] r1627_out;
	wire [31:0] r1628_out;
	wire [31:0] r1629_out;
	wire [31:0] r1630_out;
	wire [31:0] r1631_out;
	wire [31:0] r1632_out;
	wire [31:0] r1633_out;
	wire [31:0] r1634_out;
	wire [31:0] r1635_out;
	wire [31:0] r1636_out;
	wire [31:0] r1637_out;
	wire [31:0] r1638_out;
	wire [31:0] r1639_out;
	wire [31:0] r1640_out;
	wire [31:0] r1641_out;
	wire [31:0] r1642_out;
	wire [31:0] r1643_out;
	wire [31:0] r1644_out;
	wire [31:0] r1645_out;
	wire [31:0] r1646_out;
	wire [31:0] r1647_out;
	wire [31:0] r1648_out;
	wire [31:0] r1649_out;
	wire [31:0] r1650_out;
	wire [31:0] r1651_out;
	wire [31:0] r1652_out;
	wire [31:0] r1653_out;
	wire [31:0] r1654_out;
	wire [31:0] r1655_out;
	wire [31:0] r1656_out;
	wire [31:0] r1657_out;
	wire [31:0] r1658_out;
	wire [31:0] r1659_out;
	wire [31:0] r1660_out;
	wire [31:0] r1661_out;
	wire [31:0] r1662_out;
	wire [31:0] r1663_out;
	wire [31:0] r1664_out;
	wire [31:0] r1665_out;
	wire [31:0] r1666_out;
	wire [31:0] r1667_out;
	wire [31:0] r1668_out;
	wire [31:0] r1669_out;
	wire [31:0] r1670_out;
	wire [31:0] r1671_out;
	wire [31:0] r1672_out;
	wire [31:0] r1673_out;
	wire [31:0] r1674_out;
	wire [31:0] r1675_out;
	wire [31:0] r1676_out;
	wire [31:0] r1677_out;
	wire [31:0] r1678_out;
	wire [31:0] r1679_out;
	wire [31:0] r1680_out;
	wire [31:0] r1681_out;
	wire [31:0] r1682_out;
	wire [31:0] r1683_out;
	wire [31:0] r1684_out;
	wire [31:0] r1685_out;
	wire [31:0] r1686_out;
	wire [31:0] r1687_out;
	wire [31:0] r1688_out;
	wire [31:0] r1689_out;
	wire [31:0] r1690_out;
	wire [31:0] r1691_out;
	wire [31:0] r1692_out;
	wire [31:0] r1693_out;
	wire [31:0] r1694_out;
	wire [31:0] r1695_out;
	wire [31:0] r1696_out;
	wire [31:0] r1697_out;
	wire [31:0] r1698_out;
	wire [31:0] r1699_out;
	wire [31:0] r1700_out;
	wire [31:0] r1701_out;
	wire [31:0] r1702_out;
	wire [31:0] r1703_out;
	wire [31:0] r1704_out;
	wire [31:0] r1705_out;
	wire [31:0] r1706_out;
	wire [31:0] r1707_out;
	wire [31:0] r1708_out;
	wire [31:0] r1709_out;
	wire [31:0] r1710_out;
	wire [31:0] r1711_out;
	wire [31:0] r1712_out;
	wire [31:0] r1713_out;
	wire [31:0] r1714_out;
	wire [31:0] r1715_out;
	wire [31:0] r1716_out;
	wire [31:0] r1717_out;
	wire [31:0] r1718_out;
	wire [31:0] r1719_out;
	wire [31:0] r1720_out;
	wire [31:0] r1721_out;
	wire [31:0] r1722_out;
	wire [31:0] r1723_out;
	wire [31:0] r1724_out;
	wire [31:0] r1725_out;
	wire [31:0] r1726_out;
	wire [31:0] r1727_out;
	wire [31:0] r1728_out;
	wire [31:0] r1729_out;
	wire [31:0] r1730_out;
	wire [31:0] r1731_out;
	wire [31:0] r1732_out;
	wire [31:0] r1733_out;
	wire [31:0] r1734_out;
	wire [31:0] r1735_out;
	wire [31:0] r1736_out;
	wire [31:0] r1737_out;
	wire [31:0] r1738_out;
	wire [31:0] r1739_out;
	wire [31:0] r1740_out;
	wire [31:0] r1741_out;
	wire [31:0] r1742_out;
	wire [31:0] r1743_out;
	wire [31:0] r1744_out;
	wire [31:0] r1745_out;
	wire [31:0] r1746_out;
	wire [31:0] r1747_out;
	wire [31:0] r1748_out;
	wire [31:0] r1749_out;
	wire [31:0] r1750_out;
	wire [31:0] r1751_out;
	wire [31:0] r1752_out;
	wire [31:0] r1753_out;
	wire [31:0] r1754_out;
	wire [31:0] r1755_out;
	wire [31:0] r1756_out;
	wire [31:0] r1757_out;
	wire [31:0] r1758_out;
	wire [31:0] r1759_out;
	wire [31:0] r1760_out;
	wire [31:0] r1761_out;
	wire [31:0] r1762_out;
	wire [31:0] r1763_out;
	wire [31:0] r1764_out;
	wire [31:0] r1765_out;
	wire [31:0] r1766_out;
	wire [31:0] r1767_out;
	wire [31:0] r1768_out;
	wire [31:0] r1769_out;
	wire [31:0] r1770_out;
	wire [31:0] r1771_out;
	wire [31:0] r1772_out;
	wire [31:0] r1773_out;
	wire [31:0] r1774_out;
	wire [31:0] r1775_out;
	wire [31:0] r1776_out;
	wire [31:0] r1777_out;
	wire [31:0] r1778_out;
	wire [31:0] r1779_out;
	wire [31:0] r1780_out;
	wire [31:0] r1781_out;
	wire [31:0] r1782_out;
	wire [31:0] r1783_out;
	wire [31:0] r1784_out;
	wire [31:0] r1785_out;
	wire [31:0] r1786_out;
	wire [31:0] r1787_out;
	wire [31:0] r1788_out;
	wire [31:0] r1789_out;
	wire [31:0] r1790_out;
	wire [31:0] r1791_out;
	wire [31:0] r1792_out;
	wire [31:0] r1793_out;
	wire [31:0] r1794_out;
	wire [31:0] r1795_out;
	wire [31:0] r1796_out;
	wire [31:0] r1797_out;
	wire [31:0] r1798_out;
	wire [31:0] r1799_out;
	wire [31:0] r1800_out;
	wire [31:0] r1801_out;
	wire [31:0] r1802_out;
	wire [31:0] r1803_out;
	wire [31:0] r1804_out;
	wire [31:0] r1805_out;
	wire [31:0] r1806_out;
	wire [31:0] r1807_out;
	wire [31:0] r1808_out;
	wire [31:0] r1809_out;
	wire [31:0] r1810_out;
	wire [31:0] r1811_out;
	wire [31:0] r1812_out;
	wire [31:0] r1813_out;
	wire [31:0] r1814_out;
	wire [31:0] r1815_out;
	wire [31:0] r1816_out;
	wire [31:0] r1817_out;
	wire [31:0] r1818_out;
	wire [31:0] r1819_out;
	wire [31:0] r1820_out;
	wire [31:0] r1821_out;
	wire [31:0] r1822_out;
	wire [31:0] r1823_out;
	wire [31:0] r1824_out;
	wire [31:0] r1825_out;
	wire [31:0] r1826_out;
	wire [31:0] r1827_out;
	wire [31:0] r1828_out;
	wire [31:0] r1829_out;
	wire [31:0] r1830_out;
	wire [31:0] r1831_out;
	wire [31:0] r1832_out;
	wire [31:0] r1833_out;
	wire [31:0] r1834_out;
	wire [31:0] r1835_out;
	wire [31:0] r1836_out;
	wire [31:0] r1837_out;
	wire [31:0] r1838_out;
	wire [31:0] r1839_out;
	wire [31:0] r1840_out;
	wire [31:0] r1841_out;
	wire [31:0] r1842_out;
	wire [31:0] r1843_out;
	wire [31:0] r1844_out;
	wire [31:0] r1845_out;
	wire [31:0] r1846_out;
	wire [31:0] r1847_out;
	wire [31:0] r1848_out;
	wire [31:0] r1849_out;
	wire [31:0] r1850_out;
	wire [31:0] r1851_out;
	wire [31:0] r1852_out;
	wire [31:0] r1853_out;
	wire [31:0] r1854_out;
	wire [31:0] r1855_out;
	wire [31:0] r1856_out;
	wire [31:0] r1857_out;
	wire [31:0] r1858_out;
	wire [31:0] r1859_out;
	wire [31:0] r1860_out;
	wire [31:0] r1861_out;
	wire [31:0] r1862_out;
	wire [31:0] r1863_out;
	wire [31:0] r1864_out;
	wire [31:0] r1865_out;
	wire [31:0] r1866_out;
	wire [31:0] r1867_out;
	wire [31:0] r1868_out;
	wire [31:0] r1869_out;
	wire [31:0] r1870_out;
	wire [31:0] r1871_out;
	wire [31:0] r1872_out;
	wire [31:0] r1873_out;
	wire [31:0] r1874_out;
	wire [31:0] r1875_out;
	wire [31:0] r1876_out;
	wire [31:0] r1877_out;
	wire [31:0] r1878_out;
	wire [31:0] r1879_out;
	wire [31:0] r1880_out;
	wire [31:0] r1881_out;
	wire [31:0] r1882_out;
	wire [31:0] r1883_out;
	wire [31:0] r1884_out;
	wire [31:0] r1885_out;
	wire [31:0] r1886_out;
	wire [31:0] r1887_out;
	wire [31:0] r1888_out;
	wire [31:0] r1889_out;
	wire [31:0] r1890_out;
	wire [31:0] r1891_out;
	wire [31:0] r1892_out;
	wire [31:0] r1893_out;
	wire [31:0] r1894_out;
	wire [31:0] r1895_out;
	wire [31:0] r1896_out;
	wire [31:0] r1897_out;
	wire [31:0] r1898_out;
	wire [31:0] r1899_out;
	wire [31:0] r1900_out;
	wire [31:0] r1901_out;
	wire [31:0] r1902_out;
	wire [31:0] r1903_out;
	wire [31:0] r1904_out;
	wire [31:0] r1905_out;
	wire [31:0] r1906_out;
	wire [31:0] r1907_out;
	wire [31:0] r1908_out;
	wire [31:0] r1909_out;
	wire [31:0] r1910_out;
	wire [31:0] r1911_out;
	wire [31:0] r1912_out;
	wire [31:0] r1913_out;
	wire [31:0] r1914_out;
	wire [31:0] r1915_out;
	wire [31:0] r1916_out;
	wire [31:0] r1917_out;
	wire [31:0] r1918_out;
	wire [31:0] r1919_out;
	wire [31:0] r1920_out;
	wire [31:0] r1921_out;
	wire [31:0] r1922_out;
	wire [31:0] r1923_out;
	wire [31:0] r1924_out;
	wire [31:0] r1925_out;
	wire [31:0] r1926_out;
	wire [31:0] r1927_out;
	wire [31:0] r1928_out;
	wire [31:0] r1929_out;
	wire [31:0] r1930_out;
	wire [31:0] r1931_out;
	wire [31:0] r1932_out;
	wire [31:0] r1933_out;
	wire [31:0] r1934_out;
	wire [31:0] r1935_out;
	wire [31:0] r1936_out;
	wire [31:0] r1937_out;
	wire [31:0] r1938_out;
	wire [31:0] r1939_out;
	wire [31:0] r1940_out;
	wire [31:0] r1941_out;
	wire [31:0] r1942_out;
	wire [31:0] r1943_out;
	wire [31:0] r1944_out;
	wire [31:0] r1945_out;
	wire [31:0] r1946_out;
	wire [31:0] r1947_out;
	wire [31:0] r1948_out;
	wire [31:0] r1949_out;
	wire [31:0] r1950_out;
	wire [31:0] r1951_out;
	wire [31:0] r1952_out;
	wire [31:0] r1953_out;
	wire [31:0] r1954_out;
	wire [31:0] r1955_out;
	wire [31:0] r1956_out;
	wire [31:0] r1957_out;
	wire [31:0] r1958_out;
	wire [31:0] r1959_out;
	wire [31:0] r1960_out;
	wire [31:0] r1961_out;
	wire [31:0] r1962_out;
	wire [31:0] r1963_out;
	wire [31:0] r1964_out;
	wire [31:0] r1965_out;
	wire [31:0] r1966_out;
	wire [31:0] r1967_out;
	wire [31:0] r1968_out;
	wire [31:0] r1969_out;
	wire [31:0] r1970_out;
	wire [31:0] r1971_out;
	wire [31:0] r1972_out;
	wire [31:0] r1973_out;
	wire [31:0] r1974_out;
	wire [31:0] r1975_out;
	wire [31:0] r1976_out;
	wire [31:0] r1977_out;
	wire [31:0] r1978_out;
	wire [31:0] r1979_out;
	wire [31:0] r1980_out;
	wire [31:0] r1981_out;
	wire [31:0] r1982_out;
	wire [31:0] r1983_out;
	wire [31:0] r1984_out;
	wire [31:0] r1985_out;
	wire [31:0] r1986_out;
	wire [31:0] r1987_out;
	wire [31:0] r1988_out;
	wire [31:0] r1989_out;
	wire [31:0] r1990_out;
	wire [31:0] r1991_out;
	wire [31:0] r1992_out;
	wire [31:0] r1993_out;
	wire [31:0] r1994_out;
	wire [31:0] r1995_out;
	wire [31:0] r1996_out;
	wire [31:0] r1997_out;
	wire [31:0] r1998_out;
	wire [31:0] r1999_out;
	wire [31:0] r2000_out;
	wire [31:0] r2001_out;
	wire [31:0] r2002_out;
	wire [31:0] r2003_out;
	wire [31:0] r2004_out;
	wire [31:0] r2005_out;
	wire [31:0] r2006_out;
	wire [31:0] r2007_out;
	wire [31:0] r2008_out;
	wire [31:0] r2009_out;
	wire [31:0] r2010_out;
	wire [31:0] r2011_out;
	wire [31:0] r2012_out;
	wire [31:0] r2013_out;
	wire [31:0] r2014_out;
	wire [31:0] r2015_out;
	wire [31:0] r2016_out;
	wire [31:0] r2017_out;
	wire [31:0] r2018_out;
	wire [31:0] r2019_out;
	wire [31:0] r2020_out;
	wire [31:0] r2021_out;
	wire [31:0] r2022_out;
	wire [31:0] r2023_out;
	wire [31:0] r2024_out;
	wire [31:0] r2025_out;
	wire [31:0] r2026_out;
	wire [31:0] r2027_out;
	wire [31:0] r2028_out;
	wire [31:0] r2029_out;
	wire [31:0] r2030_out;
	wire [31:0] r2031_out;
	wire [31:0] r2032_out;
	wire [31:0] r2033_out;
	wire [31:0] r2034_out;
	wire [31:0] r2035_out;
	wire [31:0] r2036_out;
	wire [31:0] r2037_out;
	wire [31:0] r2038_out;
	wire [31:0] r2039_out;
	wire [31:0] r2040_out;
	wire [31:0] r2041_out;
	wire [31:0] r2042_out;
	wire [31:0] r2043_out;
	wire [31:0] r2044_out;
	wire [31:0] r2045_out;
	wire [31:0] r2046_out;
	wire [31:0] r2047_out;
	wire [31:0] r2048_out;
	wire [31:0] r2049_out;
	wire [31:0] r2050_out;
	wire [31:0] r2051_out;
	wire [31:0] r2052_out;
	wire [31:0] r2053_out;
	wire [31:0] r2054_out;
	wire [31:0] r2055_out;
	wire [31:0] r2056_out;
	wire [31:0] r2057_out;
	wire [31:0] r2058_out;
	wire [31:0] r2059_out;
	wire [31:0] r2060_out;
	wire [31:0] r2061_out;
	wire [31:0] r2062_out;
	wire [31:0] r2063_out;
	wire [31:0] r2064_out;
	wire [31:0] r2065_out;
	wire [31:0] r2066_out;
	wire [31:0] r2067_out;
	wire [31:0] r2068_out;
	wire [31:0] r2069_out;
	wire [31:0] r2070_out;
	wire [31:0] r2071_out;
	wire [31:0] r2072_out;
	wire [31:0] r2073_out;
	wire [31:0] r2074_out;
	wire [31:0] r2075_out;
	wire [31:0] r2076_out;
	wire [31:0] r2077_out;
	wire [31:0] r2078_out;
	wire [31:0] r2079_out;
	wire [31:0] r2080_out;
	wire [31:0] r2081_out;
	wire [31:0] r2082_out;
	wire [31:0] r2083_out;
	wire [31:0] r2084_out;
	wire [31:0] r2085_out;
	wire [31:0] r2086_out;
	wire [31:0] r2087_out;
	wire [31:0] r2088_out;
	wire [31:0] r2089_out;
	wire [31:0] r2090_out;
	wire [31:0] r2091_out;
	wire [31:0] r2092_out;
	wire [31:0] r2093_out;
	wire [31:0] r2094_out;
	wire [31:0] r2095_out;
	wire [31:0] r2096_out;
	wire [31:0] r2097_out;
	wire [31:0] r2098_out;
	wire [31:0] r2099_out;
	wire [31:0] r2100_out;
	wire [31:0] r2101_out;
	wire [31:0] r2102_out;
	wire [31:0] r2103_out;
	wire [31:0] r2104_out;
	wire [31:0] r2105_out;
	wire [31:0] r2106_out;
	wire [31:0] r2107_out;
	wire [31:0] r2108_out;
	wire [31:0] r2109_out;
	wire [31:0] r2110_out;
	wire [31:0] r2111_out;
	wire [31:0] r2112_out;
	wire [31:0] r2113_out;
	wire [31:0] r2114_out;
	wire [31:0] r2115_out;
	wire [31:0] r2116_out;
	wire [31:0] r2117_out;
	wire [31:0] r2118_out;
	wire [31:0] r2119_out;
	wire [31:0] r2120_out;
	wire [31:0] r2121_out;
	wire [31:0] r2122_out;
	wire [31:0] r2123_out;
	wire [31:0] r2124_out;
	wire [31:0] r2125_out;
	wire [31:0] r2126_out;
	wire [31:0] r2127_out;
	wire [31:0] r2128_out;
	wire [31:0] r2129_out;
	wire [31:0] r2130_out;
	wire [31:0] r2131_out;
	wire [31:0] r2132_out;
	wire [31:0] r2133_out;
	wire [31:0] r2134_out;
	wire [31:0] r2135_out;
	wire [31:0] r2136_out;
	wire [31:0] r2137_out;
	wire [31:0] r2138_out;
	wire [31:0] r2139_out;
	wire [31:0] r2140_out;
	wire [31:0] r2141_out;
	wire [31:0] r2142_out;
	wire [31:0] r2143_out;
	wire [31:0] r2144_out;
	wire [31:0] r2145_out;
	wire [31:0] r2146_out;
	wire [31:0] r2147_out;
	wire [31:0] r2148_out;
	wire [31:0] r2149_out;
	wire [31:0] r2150_out;
	wire [31:0] r2151_out;
	wire [31:0] r2152_out;
	wire [31:0] r2153_out;
	wire [31:0] r2154_out;
	wire [31:0] r2155_out;
	wire [31:0] r2156_out;
	wire [31:0] r2157_out;
	wire [31:0] r2158_out;
	wire [31:0] r2159_out;
	wire [31:0] r2160_out;
	wire [31:0] r2161_out;
	wire [31:0] r2162_out;
	wire [31:0] r2163_out;
	wire [31:0] r2164_out;
	wire [31:0] r2165_out;
	wire [31:0] r2166_out;
	wire [31:0] r2167_out;
	wire [31:0] r2168_out;
	wire [31:0] r2169_out;
	wire [31:0] r2170_out;
	wire [31:0] r2171_out;
	wire [31:0] r2172_out;
	wire [31:0] r2173_out;
	wire [31:0] r2174_out;
	wire [31:0] r2175_out;
	wire [31:0] r2176_out;
	wire [31:0] r2177_out;
	wire [31:0] r2178_out;
	wire [31:0] r2179_out;
	wire [31:0] r2180_out;
	wire [31:0] r2181_out;
	wire [31:0] r2182_out;
	wire [31:0] r2183_out;
	wire [31:0] r2184_out;
	wire [31:0] r2185_out;
	wire [31:0] r2186_out;
	wire [31:0] r2187_out;
	wire [31:0] r2188_out;
	wire [31:0] r2189_out;
	wire [31:0] r2190_out;
	wire [31:0] r2191_out;
	wire [31:0] r2192_out;
	wire [31:0] r2193_out;
	wire [31:0] r2194_out;
	wire [31:0] r2195_out;
	wire [31:0] r2196_out;
	wire [31:0] r2197_out;
	wire [31:0] r2198_out;
	wire [31:0] r2199_out;
	wire [31:0] r2200_out;
	wire [31:0] r2201_out;
	wire [31:0] r2202_out;
	wire [31:0] r2203_out;
	wire [31:0] r2204_out;
	wire [31:0] r2205_out;
	wire [31:0] r2206_out;
	wire [31:0] r2207_out;
	wire [31:0] r2208_out;
	wire [31:0] r2209_out;
	wire [31:0] r2210_out;
	wire [31:0] r2211_out;
	wire [31:0] r2212_out;
	wire [31:0] r2213_out;
	wire [31:0] r2214_out;
	wire [31:0] r2215_out;
	wire [31:0] r2216_out;
	wire [31:0] r2217_out;
	wire [31:0] r2218_out;
	wire [31:0] r2219_out;
	wire [31:0] r2220_out;
	wire [31:0] r2221_out;
	wire [31:0] r2222_out;
	wire [31:0] r2223_out;
	wire [31:0] r2224_out;
	wire [31:0] r2225_out;
	wire [31:0] r2226_out;
	wire [31:0] r2227_out;
	wire [31:0] r2228_out;
	wire [31:0] r2229_out;
	wire [31:0] r2230_out;
	wire [31:0] r2231_out;
	wire [31:0] r2232_out;
	wire [31:0] r2233_out;
	wire [31:0] r2234_out;
	wire [31:0] r2235_out;
	wire [31:0] r2236_out;
	wire [31:0] r2237_out;
	wire [31:0] r2238_out;
	wire [31:0] r2239_out;
	wire [31:0] r2240_out;
	wire [31:0] r2241_out;
	wire [31:0] r2242_out;
	wire [31:0] r2243_out;
	wire [31:0] r2244_out;
	wire [31:0] r2245_out;
	wire [31:0] r2246_out;
	wire [31:0] r2247_out;
	wire [31:0] r2248_out;
	wire [31:0] r2249_out;
	wire [31:0] r2250_out;
	wire [31:0] r2251_out;
	wire [31:0] r2252_out;
	wire [31:0] r2253_out;
	wire [31:0] r2254_out;
	wire [31:0] r2255_out;
	wire [31:0] r2256_out;
	wire [31:0] r2257_out;
	wire [31:0] r2258_out;
	wire [31:0] r2259_out;
	wire [31:0] r2260_out;
	wire [31:0] r2261_out;
	wire [31:0] r2262_out;
	wire [31:0] r2263_out;
	wire [31:0] r2264_out;
	wire [31:0] r2265_out;
	wire [31:0] r2266_out;
	wire [31:0] r2267_out;
	wire [31:0] r2268_out;
	wire [31:0] r2269_out;
	wire [31:0] r2270_out;
	wire [31:0] r2271_out;
	wire [31:0] r2272_out;
	wire [31:0] r2273_out;
	wire [31:0] r2274_out;
	wire [31:0] r2275_out;
	wire [31:0] r2276_out;
	wire [31:0] r2277_out;
	wire [31:0] r2278_out;
	wire [31:0] r2279_out;
	wire [31:0] r2280_out;
	wire [31:0] r2281_out;
	wire [31:0] r2282_out;
	wire [31:0] r2283_out;
	wire [31:0] r2284_out;
	wire [31:0] r2285_out;
	wire [31:0] r2286_out;
	wire [31:0] r2287_out;
	wire [31:0] r2288_out;
	wire [31:0] r2289_out;
	wire [31:0] r2290_out;
	wire [31:0] r2291_out;
	wire [31:0] r2292_out;
	wire [31:0] r2293_out;
	wire [31:0] r2294_out;
	wire [31:0] r2295_out;
	wire [31:0] r2296_out;
	wire [31:0] r2297_out;
	wire [31:0] r2298_out;
	wire [31:0] r2299_out;
	wire [31:0] r2300_out;
	wire [31:0] r2301_out;
	wire [31:0] r2302_out;
	wire [31:0] r2303_out;
	wire [31:0] r2304_out;
	wire [31:0] r2305_out;
	wire [31:0] r2306_out;
	wire [31:0] r2307_out;
	wire [31:0] r2308_out;
	wire [31:0] r2309_out;
	wire [31:0] r2310_out;
	wire [31:0] r2311_out;
	wire [31:0] r2312_out;
	wire [31:0] r2313_out;
	wire [31:0] r2314_out;
	wire [31:0] r2315_out;
	wire [31:0] r2316_out;
	wire [31:0] r2317_out;
	wire [31:0] r2318_out;
	wire [31:0] r2319_out;
	wire [31:0] r2320_out;
	wire [31:0] r2321_out;
	wire [31:0] r2322_out;
	wire [31:0] r2323_out;
	wire [31:0] r2324_out;
	wire [31:0] r2325_out;
	wire [31:0] r2326_out;
	wire [31:0] r2327_out;
	wire [31:0] r2328_out;
	wire [31:0] r2329_out;
	wire [31:0] r2330_out;
	wire [31:0] r2331_out;
	wire [31:0] r2332_out;
	wire [31:0] r2333_out;
	wire [31:0] r2334_out;
	wire [31:0] r2335_out;
	wire [31:0] r2336_out;
	wire [31:0] r2337_out;
	wire [31:0] r2338_out;
	wire [31:0] r2339_out;
	wire [31:0] r2340_out;
	wire [31:0] r2341_out;
	wire [31:0] r2342_out;
	wire [31:0] r2343_out;
	wire [31:0] r2344_out;
	wire [31:0] r2345_out;
	wire [31:0] r2346_out;
	wire [31:0] r2347_out;
	wire [31:0] r2348_out;
	wire [31:0] r2349_out;
	wire [31:0] r2350_out;
	wire [31:0] r2351_out;
	wire [31:0] r2352_out;
	wire [31:0] r2353_out;
	wire [31:0] r2354_out;
	wire [31:0] r2355_out;
	wire [31:0] r2356_out;
	wire [31:0] r2357_out;
	wire [31:0] r2358_out;
	wire [31:0] r2359_out;
	wire [31:0] r2360_out;
	wire [31:0] r2361_out;
	wire [31:0] r2362_out;
	wire [31:0] r2363_out;
	wire [31:0] r2364_out;
	wire [31:0] r2365_out;
	wire [31:0] r2366_out;
	wire [31:0] r2367_out;
	wire [31:0] r2368_out;
	wire [31:0] r2369_out;
	wire [31:0] r2370_out;
	wire [31:0] r2371_out;
	wire [31:0] r2372_out;
	wire [31:0] r2373_out;
	wire [31:0] r2374_out;
	wire [31:0] r2375_out;
	wire [31:0] r2376_out;
	wire [31:0] r2377_out;
	wire [31:0] r2378_out;
	wire [31:0] r2379_out;
	wire [31:0] r2380_out;
	wire [31:0] r2381_out;
	wire [31:0] r2382_out;
	wire [31:0] r2383_out;
	wire [31:0] r2384_out;
	wire [31:0] r2385_out;
	wire [31:0] r2386_out;
	wire [31:0] r2387_out;
	wire [31:0] r2388_out;
	wire [31:0] r2389_out;
	wire [31:0] r2390_out;
	wire [31:0] r2391_out;
	wire [31:0] r2392_out;
	wire [31:0] r2393_out;
	wire [31:0] r2394_out;
	wire [31:0] r2395_out;
	wire [31:0] r2396_out;
	wire [31:0] r2397_out;
	wire [31:0] r2398_out;
	wire [31:0] r2399_out;
	wire [31:0] r2400_out;
	wire [31:0] r2401_out;
	wire [31:0] r2402_out;
	wire [31:0] r2403_out;
	wire [31:0] r2404_out;
	wire [31:0] r2405_out;
	wire [31:0] r2406_out;
	wire [31:0] r2407_out;
	wire [31:0] r2408_out;
	wire [31:0] r2409_out;
	wire [31:0] r2410_out;
	wire [31:0] r2411_out;
	wire [31:0] r2412_out;
	wire [31:0] r2413_out;
	wire [31:0] r2414_out;
	wire [31:0] r2415_out;
	wire [31:0] r2416_out;
	wire [31:0] r2417_out;
	wire [31:0] r2418_out;
	wire [31:0] r2419_out;
	wire [31:0] r2420_out;
	wire [31:0] r2421_out;
	wire [31:0] r2422_out;
	wire [31:0] r2423_out;
	wire [31:0] r2424_out;
	wire [31:0] r2425_out;
	wire [31:0] r2426_out;
	wire [31:0] r2427_out;
	wire [31:0] r2428_out;
	wire [31:0] r2429_out;
	wire [31:0] r2430_out;
	wire [31:0] r2431_out;
	wire [31:0] r2432_out;
	wire [31:0] r2433_out;
	wire [31:0] r2434_out;
	wire [31:0] r2435_out;
	wire [31:0] r2436_out;
	wire [31:0] r2437_out;
	wire [31:0] r2438_out;
	wire [31:0] r2439_out;
	wire [31:0] r2440_out;
	wire [31:0] r2441_out;
	wire [31:0] r2442_out;
	wire [31:0] r2443_out;
	wire [31:0] r2444_out;
	wire [31:0] r2445_out;
	wire [31:0] r2446_out;
	wire [31:0] r2447_out;
	wire [31:0] r2448_out;
	wire [31:0] r2449_out;
	wire [31:0] r2450_out;
	wire [31:0] r2451_out;
	wire [31:0] r2452_out;
	wire [31:0] r2453_out;
	wire [31:0] r2454_out;
	wire [31:0] r2455_out;
	wire [31:0] r2456_out;
	wire [31:0] r2457_out;
	wire [31:0] r2458_out;
	wire [31:0] r2459_out;
	wire [31:0] r2460_out;
	wire [31:0] r2461_out;
	wire [31:0] r2462_out;
	wire [31:0] r2463_out;
	wire [31:0] r2464_out;
	wire [31:0] r2465_out;
	wire [31:0] r2466_out;
	wire [31:0] r2467_out;
	wire [31:0] r2468_out;
	wire [31:0] r2469_out;
	wire [31:0] r2470_out;
	wire [31:0] r2471_out;
	wire [31:0] r2472_out;
	wire [31:0] r2473_out;
	wire [31:0] r2474_out;
	wire [31:0] r2475_out;
	wire [31:0] r2476_out;
	wire [31:0] r2477_out;
	wire [31:0] r2478_out;
	wire [31:0] r2479_out;
	wire [31:0] r2480_out;
	wire [31:0] r2481_out;
	wire [31:0] r2482_out;
	wire [31:0] r2483_out;
	wire [31:0] r2484_out;
	wire [31:0] r2485_out;
	wire [31:0] r2486_out;
	wire [31:0] r2487_out;
	wire [31:0] r2488_out;
	wire [31:0] r2489_out;
	wire [31:0] r2490_out;
	wire [31:0] r2491_out;
	wire [31:0] r2492_out;
	wire [31:0] r2493_out;
	wire [31:0] r2494_out;
	wire [31:0] r2495_out;
	wire [31:0] r2496_out;
	wire [31:0] r2497_out;
	wire [31:0] r2498_out;
	wire [31:0] r2499_out;
	wire [31:0] r2500_out;
	wire [31:0] r2501_out;
	wire [31:0] r2502_out;
	wire [31:0] r2503_out;
	wire [31:0] r2504_out;
	wire [31:0] r2505_out;
	wire [31:0] r2506_out;
	wire [31:0] r2507_out;
	wire [31:0] r2508_out;
	wire [31:0] r2509_out;
	wire [31:0] r2510_out;
	wire [31:0] r2511_out;
	wire [31:0] r2512_out;
	wire [31:0] r2513_out;
	wire [31:0] r2514_out;
	wire [31:0] r2515_out;
	wire [31:0] r2516_out;
	wire [31:0] r2517_out;
	wire [31:0] r2518_out;
	wire [31:0] r2519_out;
	wire [31:0] r2520_out;
	wire [31:0] r2521_out;
	wire [31:0] r2522_out;
	wire [31:0] r2523_out;
	wire [31:0] r2524_out;
	wire [31:0] r2525_out;
	wire [31:0] r2526_out;
	wire [31:0] r2527_out;
	wire [31:0] r2528_out;
	wire [31:0] r2529_out;
	wire [31:0] r2530_out;
	wire [31:0] r2531_out;
	wire [31:0] r2532_out;
	wire [31:0] r2533_out;
	wire [31:0] r2534_out;
	wire [31:0] r2535_out;
	wire [31:0] r2536_out;
	wire [31:0] r2537_out;
	wire [31:0] r2538_out;
	wire [31:0] r2539_out;
	wire [31:0] r2540_out;
	wire [31:0] r2541_out;
	wire [31:0] r2542_out;
	wire [31:0] r2543_out;
	wire [31:0] r2544_out;
	wire [31:0] r2545_out;
	wire [31:0] r2546_out;
	wire [31:0] r2547_out;
	wire [31:0] r2548_out;
	wire [31:0] r2549_out;
	wire [31:0] r2550_out;
	wire [31:0] r2551_out;
	wire [31:0] r2552_out;
	wire [31:0] r2553_out;
	wire [31:0] r2554_out;
	wire [31:0] r2555_out;
	wire [31:0] r2556_out;
	wire [31:0] r2557_out;
	wire [31:0] r2558_out;
	wire [31:0] r2559_out;
	wire [31:0] r2560_out;
	wire [31:0] r2561_out;
	wire [31:0] r2562_out;
	wire [31:0] r2563_out;
	wire [31:0] r2564_out;
	wire [31:0] r2565_out;
	wire [31:0] r2566_out;
	wire [31:0] r2567_out;
	wire [31:0] r2568_out;
	wire [31:0] r2569_out;
	wire [31:0] r2570_out;
	wire [31:0] r2571_out;
	wire [31:0] r2572_out;
	wire [31:0] r2573_out;
	wire [31:0] r2574_out;
	wire [31:0] r2575_out;
	wire [31:0] r2576_out;
	wire [31:0] r2577_out;
	wire [31:0] r2578_out;
	wire [31:0] r2579_out;
	wire [31:0] r2580_out;
	wire [31:0] r2581_out;
	wire [31:0] r2582_out;
	wire [31:0] r2583_out;
	wire [31:0] r2584_out;
	wire [31:0] r2585_out;
	wire [31:0] r2586_out;
	wire [31:0] r2587_out;
	wire [31:0] r2588_out;
	wire [31:0] r2589_out;
	wire [31:0] r2590_out;
	wire [31:0] r2591_out;
	wire [31:0] r2592_out;
	wire [31:0] r2593_out;
	wire [31:0] r2594_out;
	wire [31:0] r2595_out;
	wire [31:0] r2596_out;
	wire [31:0] r2597_out;
	wire [31:0] r2598_out;
	wire [31:0] r2599_out;
	wire [31:0] r2600_out;
	wire [31:0] r2601_out;
	wire [31:0] r2602_out;
	wire [31:0] r2603_out;
	wire [31:0] r2604_out;
	wire [31:0] r2605_out;
	wire [31:0] r2606_out;
	wire [31:0] r2607_out;
	wire [31:0] r2608_out;
	wire [31:0] r2609_out;
	wire [31:0] r2610_out;
	wire [31:0] r2611_out;
	wire [31:0] r2612_out;
	wire [31:0] r2613_out;
	wire [31:0] r2614_out;
	wire [31:0] r2615_out;
	wire [31:0] r2616_out;
	wire [31:0] r2617_out;
	wire [31:0] r2618_out;
	wire [31:0] r2619_out;
	wire [31:0] r2620_out;
	wire [31:0] r2621_out;
	wire [31:0] r2622_out;
	wire [31:0] r2623_out;
	wire [31:0] r2624_out;
	wire [31:0] r2625_out;
	wire [31:0] r2626_out;
	wire [31:0] r2627_out;
	wire [31:0] r2628_out;
	wire [31:0] r2629_out;
	wire [31:0] r2630_out;
	wire [31:0] r2631_out;
	wire [31:0] r2632_out;
	wire [31:0] r2633_out;
	wire [31:0] r2634_out;
	wire [31:0] r2635_out;
	wire [31:0] r2636_out;
	wire [31:0] r2637_out;
	wire [31:0] r2638_out;
	wire [31:0] r2639_out;
	wire [31:0] r2640_out;
	wire [31:0] r2641_out;
	wire [31:0] r2642_out;
	wire [31:0] r2643_out;
	wire [31:0] r2644_out;
	wire [31:0] r2645_out;
	wire [31:0] r2646_out;
	wire [31:0] r2647_out;
	wire [31:0] r2648_out;
	wire [31:0] r2649_out;
	wire [31:0] r2650_out;
	wire [31:0] r2651_out;
	wire [31:0] r2652_out;
	wire [31:0] r2653_out;
	wire [31:0] r2654_out;
	wire [31:0] r2655_out;
	wire [31:0] r2656_out;
	wire [31:0] r2657_out;
	wire [31:0] r2658_out;
	wire [31:0] r2659_out;
	wire [31:0] r2660_out;
	wire [31:0] r2661_out;
	wire [31:0] r2662_out;
	wire [31:0] r2663_out;
	wire [31:0] r2664_out;
	wire [31:0] r2665_out;
	wire [31:0] r2666_out;
	wire [31:0] r2667_out;
	wire [31:0] r2668_out;
	wire [31:0] r2669_out;
	wire [31:0] r2670_out;
	wire [31:0] r2671_out;
	wire [31:0] r2672_out;
	wire [31:0] r2673_out;
	wire [31:0] r2674_out;
	wire [31:0] r2675_out;
	wire [31:0] r2676_out;
	wire [31:0] r2677_out;
	wire [31:0] r2678_out;
	wire [31:0] r2679_out;
	wire [31:0] r2680_out;
	wire [31:0] r2681_out;
	wire [31:0] r2682_out;
	wire [31:0] r2683_out;
	wire [31:0] r2684_out;
	wire [31:0] r2685_out;
	wire [31:0] r2686_out;
	wire [31:0] r2687_out;
	wire [31:0] r2688_out;
	wire [31:0] r2689_out;
	wire [31:0] r2690_out;
	wire [31:0] r2691_out;
	wire [31:0] r2692_out;
	wire [31:0] r2693_out;
	wire [31:0] r2694_out;
	wire [31:0] r2695_out;
	wire [31:0] r2696_out;
	wire [31:0] r2697_out;
	wire [31:0] r2698_out;
	wire [31:0] r2699_out;
	wire [31:0] r2700_out;
	wire [31:0] r2701_out;
	wire [31:0] r2702_out;
	wire [31:0] r2703_out;
	wire [31:0] r2704_out;
	wire [31:0] r2705_out;
	wire [31:0] r2706_out;
	wire [31:0] r2707_out;
	wire [31:0] r2708_out;
	wire [31:0] r2709_out;
	wire [31:0] r2710_out;
	wire [31:0] r2711_out;
	wire [31:0] r2712_out;
	wire [31:0] r2713_out;
	wire [31:0] r2714_out;
	wire [31:0] r2715_out;
	wire [31:0] r2716_out;
	wire [31:0] r2717_out;
	wire [31:0] r2718_out;
	wire [31:0] r2719_out;
	wire [31:0] r2720_out;
	wire [31:0] r2721_out;
	wire [31:0] r2722_out;
	wire [31:0] r2723_out;
	wire [31:0] r2724_out;
	wire [31:0] r2725_out;
	wire [31:0] r2726_out;
	wire [31:0] r2727_out;
	wire [31:0] r2728_out;
	wire [31:0] r2729_out;
	wire [31:0] r2730_out;
	wire [31:0] r2731_out;
	wire [31:0] r2732_out;
	wire [31:0] r2733_out;
	wire [31:0] r2734_out;
	wire [31:0] r2735_out;
	wire [31:0] r2736_out;
	wire [31:0] r2737_out;
	wire [31:0] r2738_out;
	wire [31:0] r2739_out;
	wire [31:0] r2740_out;
	wire [31:0] r2741_out;
	wire [31:0] r2742_out;
	wire [31:0] r2743_out;
	wire [31:0] r2744_out;
	wire [31:0] r2745_out;
	wire [31:0] r2746_out;
	wire [31:0] r2747_out;
	wire [31:0] r2748_out;
	wire [31:0] r2749_out;
	wire [31:0] r2750_out;
	wire [31:0] r2751_out;
	wire [31:0] r2752_out;
	wire [31:0] r2753_out;
	wire [31:0] r2754_out;
	wire [31:0] r2755_out;
	wire [31:0] r2756_out;
	wire [31:0] r2757_out;
	wire [31:0] r2758_out;
	wire [31:0] r2759_out;
	wire [31:0] r2760_out;
	wire [31:0] r2761_out;
	wire [31:0] r2762_out;
	wire [31:0] r2763_out;
	wire [31:0] r2764_out;
	wire [31:0] r2765_out;
	wire [31:0] r2766_out;
	wire [31:0] r2767_out;
	wire [31:0] r2768_out;
	wire [31:0] r2769_out;
	wire [31:0] r2770_out;
	wire [31:0] r2771_out;
	wire [31:0] r2772_out;
	wire [31:0] r2773_out;
	wire [31:0] r2774_out;
	wire [31:0] r2775_out;
	wire [31:0] r2776_out;
	wire [31:0] r2777_out;
	wire [31:0] r2778_out;
	wire [31:0] r2779_out;
	wire [31:0] r2780_out;
	wire [31:0] r2781_out;
	wire [31:0] r2782_out;
	wire [31:0] r2783_out;
	wire [31:0] r2784_out;
	wire [31:0] r2785_out;
	wire [31:0] r2786_out;
	wire [31:0] r2787_out;
	wire [31:0] r2788_out;
	wire [31:0] r2789_out;
	wire [31:0] r2790_out;
	wire [31:0] r2791_out;
	wire [31:0] r2792_out;
	wire [31:0] r2793_out;
	wire [31:0] r2794_out;
	wire [31:0] r2795_out;
	wire [31:0] r2796_out;
	wire [31:0] r2797_out;
	wire [31:0] r2798_out;
	wire [31:0] r2799_out;
	wire [31:0] r2800_out;
	wire [31:0] r2801_out;
	wire [31:0] r2802_out;
	wire [31:0] r2803_out;
	wire [31:0] r2804_out;
	wire [31:0] r2805_out;
	wire [31:0] r2806_out;
	wire [31:0] r2807_out;
	wire [31:0] r2808_out;
	wire [31:0] r2809_out;
	wire [31:0] r2810_out;
	wire [31:0] r2811_out;
	wire [31:0] r2812_out;
	wire [31:0] r2813_out;
	wire [31:0] r2814_out;
	wire [31:0] r2815_out;
	wire [31:0] r2816_out;
	wire [31:0] r2817_out;
	wire [31:0] r2818_out;
	wire [31:0] r2819_out;
	wire [31:0] r2820_out;
	wire [31:0] r2821_out;
	wire [31:0] r2822_out;
	wire [31:0] r2823_out;
	wire [31:0] r2824_out;
	wire [31:0] r2825_out;
	wire [31:0] r2826_out;
	wire [31:0] r2827_out;
	wire [31:0] r2828_out;
	wire [31:0] r2829_out;
	wire [31:0] r2830_out;
	wire [31:0] r2831_out;
	wire [31:0] r2832_out;
	wire [31:0] r2833_out;
	wire [31:0] r2834_out;
	wire [31:0] r2835_out;
	wire [31:0] r2836_out;
	wire [31:0] r2837_out;
	wire [31:0] r2838_out;
	wire [31:0] r2839_out;
	wire [31:0] r2840_out;
	wire [31:0] r2841_out;
	wire [31:0] r2842_out;
	wire [31:0] r2843_out;
	wire [31:0] r2844_out;
	wire [31:0] r2845_out;
	wire [31:0] r2846_out;
	wire [31:0] r2847_out;
	wire [31:0] r2848_out;
	wire [31:0] r2849_out;
	wire [31:0] r2850_out;
	wire [31:0] r2851_out;
	wire [31:0] r2852_out;
	wire [31:0] r2853_out;
	wire [31:0] r2854_out;
	wire [31:0] r2855_out;
	wire [31:0] r2856_out;
	wire [31:0] r2857_out;
	wire [31:0] r2858_out;
	wire [31:0] r2859_out;
	wire [31:0] r2860_out;
	wire [31:0] r2861_out;
	wire [31:0] r2862_out;
	wire [31:0] r2863_out;
	wire [31:0] r2864_out;
	wire [31:0] r2865_out;
	wire [31:0] r2866_out;
	wire [31:0] r2867_out;
	wire [31:0] r2868_out;
	wire [31:0] r2869_out;
	wire [31:0] r2870_out;
	wire [31:0] r2871_out;
	wire [31:0] r2872_out;
	wire [31:0] r2873_out;
	wire [31:0] r2874_out;
	wire [31:0] r2875_out;
	wire [31:0] r2876_out;
	wire [31:0] r2877_out;
	wire [31:0] r2878_out;
	wire [31:0] r2879_out;
	wire [31:0] r2880_out;
	wire [31:0] r2881_out;
	wire [31:0] r2882_out;
	wire [31:0] r2883_out;
	wire [31:0] r2884_out;
	wire [31:0] r2885_out;
	wire [31:0] r2886_out;
	wire [31:0] r2887_out;
	wire [31:0] r2888_out;
	wire [31:0] r2889_out;
	wire [31:0] r2890_out;
	wire [31:0] r2891_out;
	wire [31:0] r2892_out;
	wire [31:0] r2893_out;
	wire [31:0] r2894_out;
	wire [31:0] r2895_out;
	wire [31:0] r2896_out;
	wire [31:0] r2897_out;
	wire [31:0] r2898_out;
	wire [31:0] r2899_out;
	wire [31:0] r2900_out;
	wire [31:0] r2901_out;
	wire [31:0] r2902_out;
	wire [31:0] r2903_out;
	wire [31:0] r2904_out;
	wire [31:0] r2905_out;
	wire [31:0] r2906_out;
	wire [31:0] r2907_out;
	wire [31:0] r2908_out;
	wire [31:0] r2909_out;
	wire [31:0] r2910_out;
	wire [31:0] r2911_out;
	wire [31:0] r2912_out;
	wire [31:0] r2913_out;
	wire [31:0] r2914_out;
	wire [31:0] r2915_out;
	wire [31:0] r2916_out;
	wire [31:0] r2917_out;
	wire [31:0] r2918_out;
	wire [31:0] r2919_out;
	wire [31:0] r2920_out;
	wire [31:0] r2921_out;
	wire [31:0] r2922_out;
	wire [31:0] r2923_out;
	wire [31:0] r2924_out;
	wire [31:0] r2925_out;
	wire [31:0] r2926_out;
	wire [31:0] r2927_out;
	wire [31:0] r2928_out;
	wire [31:0] r2929_out;
	wire [31:0] r2930_out;
	wire [31:0] r2931_out;
	wire [31:0] r2932_out;
	wire [31:0] r2933_out;
	wire [31:0] r2934_out;
	wire [31:0] r2935_out;
	wire [31:0] r2936_out;
	wire [31:0] r2937_out;
	wire [31:0] r2938_out;
	wire [31:0] r2939_out;
	wire [31:0] r2940_out;
	wire [31:0] r2941_out;
	wire [31:0] r2942_out;
	wire [31:0] r2943_out;
	wire [31:0] r2944_out;
	wire [31:0] r2945_out;
	wire [31:0] r2946_out;
	wire [31:0] r2947_out;
	wire [31:0] r2948_out;
	wire [31:0] r2949_out;
	wire [31:0] r2950_out;
	wire [31:0] r2951_out;
	wire [31:0] r2952_out;
	wire [31:0] r2953_out;
	wire [31:0] r2954_out;
	wire [31:0] r2955_out;
	wire [31:0] r2956_out;
	wire [31:0] r2957_out;
	wire [31:0] r2958_out;
	wire [31:0] r2959_out;
	wire [31:0] r2960_out;
	wire [31:0] r2961_out;
	wire [31:0] r2962_out;
	wire [31:0] r2963_out;
	wire [31:0] r2964_out;
	wire [31:0] r2965_out;
	wire [31:0] r2966_out;
	wire [31:0] r2967_out;
	wire [31:0] r2968_out;
	wire [31:0] r2969_out;
	wire [31:0] r2970_out;
	wire [31:0] r2971_out;
	wire [31:0] r2972_out;
	wire [31:0] r2973_out;
	wire [31:0] r2974_out;
	wire [31:0] r2975_out;
	wire [31:0] r2976_out;
	wire [31:0] r2977_out;
	wire [31:0] r2978_out;
	wire [31:0] r2979_out;
	wire [31:0] r2980_out;
	wire [31:0] r2981_out;
	wire [31:0] r2982_out;
	wire [31:0] r2983_out;
	wire [31:0] r2984_out;
	wire [31:0] r2985_out;
	wire [31:0] r2986_out;
	wire [31:0] r2987_out;
	wire [31:0] r2988_out;
	wire [31:0] r2989_out;
	wire [31:0] r2990_out;
	wire [31:0] r2991_out;
	wire [31:0] r2992_out;
	wire [31:0] r2993_out;
	wire [31:0] r2994_out;
	wire [31:0] r2995_out;
	wire [31:0] r2996_out;
	wire [31:0] r2997_out;
	wire [31:0] r2998_out;
	wire [31:0] r2999_out;

	reg32 r0 (rst, clk, in, r0_out);
	reg32 r1 (rst, clk, r0_out, r1_out);
	reg32 r2 (rst, clk, r1_out, r2_out);
	reg32 r3 (rst, clk, r2_out, r3_out);
	reg32 r4 (rst, clk, r3_out, r4_out);
	reg32 r5 (rst, clk, r4_out, r5_out);
	reg32 r6 (rst, clk, r5_out, r6_out);
	reg32 r7 (rst, clk, r6_out, r7_out);
	reg32 r8 (rst, clk, r7_out, r8_out);
	reg32 r9 (rst, clk, r8_out, r9_out);
	reg32 r10 (rst, clk, r9_out, r10_out);
	reg32 r11 (rst, clk, r10_out, r11_out);
	reg32 r12 (rst, clk, r11_out, r12_out);
	reg32 r13 (rst, clk, r12_out, r13_out);
	reg32 r14 (rst, clk, r13_out, r14_out);
	reg32 r15 (rst, clk, r14_out, r15_out);
	reg32 r16 (rst, clk, r15_out, r16_out);
	reg32 r17 (rst, clk, r16_out, r17_out);
	reg32 r18 (rst, clk, r17_out, r18_out);
	reg32 r19 (rst, clk, r18_out, r19_out);
	reg32 r20 (rst, clk, r19_out, r20_out);
	reg32 r21 (rst, clk, r20_out, r21_out);
	reg32 r22 (rst, clk, r21_out, r22_out);
	reg32 r23 (rst, clk, r22_out, r23_out);
	reg32 r24 (rst, clk, r23_out, r24_out);
	reg32 r25 (rst, clk, r24_out, r25_out);
	reg32 r26 (rst, clk, r25_out, r26_out);
	reg32 r27 (rst, clk, r26_out, r27_out);
	reg32 r28 (rst, clk, r27_out, r28_out);
	reg32 r29 (rst, clk, r28_out, r29_out);
	reg32 r30 (rst, clk, r29_out, r30_out);
	reg32 r31 (rst, clk, r30_out, r31_out);
	reg32 r32 (rst, clk, r31_out, r32_out);
	reg32 r33 (rst, clk, r32_out, r33_out);
	reg32 r34 (rst, clk, r33_out, r34_out);
	reg32 r35 (rst, clk, r34_out, r35_out);
	reg32 r36 (rst, clk, r35_out, r36_out);
	reg32 r37 (rst, clk, r36_out, r37_out);
	reg32 r38 (rst, clk, r37_out, r38_out);
	reg32 r39 (rst, clk, r38_out, r39_out);
	reg32 r40 (rst, clk, r39_out, r40_out);
	reg32 r41 (rst, clk, r40_out, r41_out);
	reg32 r42 (rst, clk, r41_out, r42_out);
	reg32 r43 (rst, clk, r42_out, r43_out);
	reg32 r44 (rst, clk, r43_out, r44_out);
	reg32 r45 (rst, clk, r44_out, r45_out);
	reg32 r46 (rst, clk, r45_out, r46_out);
	reg32 r47 (rst, clk, r46_out, r47_out);
	reg32 r48 (rst, clk, r47_out, r48_out);
	reg32 r49 (rst, clk, r48_out, r49_out);
	reg32 r50 (rst, clk, r49_out, r50_out);
	reg32 r51 (rst, clk, r50_out, r51_out);
	reg32 r52 (rst, clk, r51_out, r52_out);
	reg32 r53 (rst, clk, r52_out, r53_out);
	reg32 r54 (rst, clk, r53_out, r54_out);
	reg32 r55 (rst, clk, r54_out, r55_out);
	reg32 r56 (rst, clk, r55_out, r56_out);
	reg32 r57 (rst, clk, r56_out, r57_out);
	reg32 r58 (rst, clk, r57_out, r58_out);
	reg32 r59 (rst, clk, r58_out, r59_out);
	reg32 r60 (rst, clk, r59_out, r60_out);
	reg32 r61 (rst, clk, r60_out, r61_out);
	reg32 r62 (rst, clk, r61_out, r62_out);
	reg32 r63 (rst, clk, r62_out, r63_out);
	reg32 r64 (rst, clk, r63_out, r64_out);
	reg32 r65 (rst, clk, r64_out, r65_out);
	reg32 r66 (rst, clk, r65_out, r66_out);
	reg32 r67 (rst, clk, r66_out, r67_out);
	reg32 r68 (rst, clk, r67_out, r68_out);
	reg32 r69 (rst, clk, r68_out, r69_out);
	reg32 r70 (rst, clk, r69_out, r70_out);
	reg32 r71 (rst, clk, r70_out, r71_out);
	reg32 r72 (rst, clk, r71_out, r72_out);
	reg32 r73 (rst, clk, r72_out, r73_out);
	reg32 r74 (rst, clk, r73_out, r74_out);
	reg32 r75 (rst, clk, r74_out, r75_out);
	reg32 r76 (rst, clk, r75_out, r76_out);
	reg32 r77 (rst, clk, r76_out, r77_out);
	reg32 r78 (rst, clk, r77_out, r78_out);
	reg32 r79 (rst, clk, r78_out, r79_out);
	reg32 r80 (rst, clk, r79_out, r80_out);
	reg32 r81 (rst, clk, r80_out, r81_out);
	reg32 r82 (rst, clk, r81_out, r82_out);
	reg32 r83 (rst, clk, r82_out, r83_out);
	reg32 r84 (rst, clk, r83_out, r84_out);
	reg32 r85 (rst, clk, r84_out, r85_out);
	reg32 r86 (rst, clk, r85_out, r86_out);
	reg32 r87 (rst, clk, r86_out, r87_out);
	reg32 r88 (rst, clk, r87_out, r88_out);
	reg32 r89 (rst, clk, r88_out, r89_out);
	reg32 r90 (rst, clk, r89_out, r90_out);
	reg32 r91 (rst, clk, r90_out, r91_out);
	reg32 r92 (rst, clk, r91_out, r92_out);
	reg32 r93 (rst, clk, r92_out, r93_out);
	reg32 r94 (rst, clk, r93_out, r94_out);
	reg32 r95 (rst, clk, r94_out, r95_out);
	reg32 r96 (rst, clk, r95_out, r96_out);
	reg32 r97 (rst, clk, r96_out, r97_out);
	reg32 r98 (rst, clk, r97_out, r98_out);
	reg32 r99 (rst, clk, r98_out, r99_out);
	reg32 r100 (rst, clk, r99_out, r100_out);
	reg32 r101 (rst, clk, r100_out, r101_out);
	reg32 r102 (rst, clk, r101_out, r102_out);
	reg32 r103 (rst, clk, r102_out, r103_out);
	reg32 r104 (rst, clk, r103_out, r104_out);
	reg32 r105 (rst, clk, r104_out, r105_out);
	reg32 r106 (rst, clk, r105_out, r106_out);
	reg32 r107 (rst, clk, r106_out, r107_out);
	reg32 r108 (rst, clk, r107_out, r108_out);
	reg32 r109 (rst, clk, r108_out, r109_out);
	reg32 r110 (rst, clk, r109_out, r110_out);
	reg32 r111 (rst, clk, r110_out, r111_out);
	reg32 r112 (rst, clk, r111_out, r112_out);
	reg32 r113 (rst, clk, r112_out, r113_out);
	reg32 r114 (rst, clk, r113_out, r114_out);
	reg32 r115 (rst, clk, r114_out, r115_out);
	reg32 r116 (rst, clk, r115_out, r116_out);
	reg32 r117 (rst, clk, r116_out, r117_out);
	reg32 r118 (rst, clk, r117_out, r118_out);
	reg32 r119 (rst, clk, r118_out, r119_out);
	reg32 r120 (rst, clk, r119_out, r120_out);
	reg32 r121 (rst, clk, r120_out, r121_out);
	reg32 r122 (rst, clk, r121_out, r122_out);
	reg32 r123 (rst, clk, r122_out, r123_out);
	reg32 r124 (rst, clk, r123_out, r124_out);
	reg32 r125 (rst, clk, r124_out, r125_out);
	reg32 r126 (rst, clk, r125_out, r126_out);
	reg32 r127 (rst, clk, r126_out, r127_out);
	reg32 r128 (rst, clk, r127_out, r128_out);
	reg32 r129 (rst, clk, r128_out, r129_out);
	reg32 r130 (rst, clk, r129_out, r130_out);
	reg32 r131 (rst, clk, r130_out, r131_out);
	reg32 r132 (rst, clk, r131_out, r132_out);
	reg32 r133 (rst, clk, r132_out, r133_out);
	reg32 r134 (rst, clk, r133_out, r134_out);
	reg32 r135 (rst, clk, r134_out, r135_out);
	reg32 r136 (rst, clk, r135_out, r136_out);
	reg32 r137 (rst, clk, r136_out, r137_out);
	reg32 r138 (rst, clk, r137_out, r138_out);
	reg32 r139 (rst, clk, r138_out, r139_out);
	reg32 r140 (rst, clk, r139_out, r140_out);
	reg32 r141 (rst, clk, r140_out, r141_out);
	reg32 r142 (rst, clk, r141_out, r142_out);
	reg32 r143 (rst, clk, r142_out, r143_out);
	reg32 r144 (rst, clk, r143_out, r144_out);
	reg32 r145 (rst, clk, r144_out, r145_out);
	reg32 r146 (rst, clk, r145_out, r146_out);
	reg32 r147 (rst, clk, r146_out, r147_out);
	reg32 r148 (rst, clk, r147_out, r148_out);
	reg32 r149 (rst, clk, r148_out, r149_out);
	reg32 r150 (rst, clk, r149_out, r150_out);
	reg32 r151 (rst, clk, r150_out, r151_out);
	reg32 r152 (rst, clk, r151_out, r152_out);
	reg32 r153 (rst, clk, r152_out, r153_out);
	reg32 r154 (rst, clk, r153_out, r154_out);
	reg32 r155 (rst, clk, r154_out, r155_out);
	reg32 r156 (rst, clk, r155_out, r156_out);
	reg32 r157 (rst, clk, r156_out, r157_out);
	reg32 r158 (rst, clk, r157_out, r158_out);
	reg32 r159 (rst, clk, r158_out, r159_out);
	reg32 r160 (rst, clk, r159_out, r160_out);
	reg32 r161 (rst, clk, r160_out, r161_out);
	reg32 r162 (rst, clk, r161_out, r162_out);
	reg32 r163 (rst, clk, r162_out, r163_out);
	reg32 r164 (rst, clk, r163_out, r164_out);
	reg32 r165 (rst, clk, r164_out, r165_out);
	reg32 r166 (rst, clk, r165_out, r166_out);
	reg32 r167 (rst, clk, r166_out, r167_out);
	reg32 r168 (rst, clk, r167_out, r168_out);
	reg32 r169 (rst, clk, r168_out, r169_out);
	reg32 r170 (rst, clk, r169_out, r170_out);
	reg32 r171 (rst, clk, r170_out, r171_out);
	reg32 r172 (rst, clk, r171_out, r172_out);
	reg32 r173 (rst, clk, r172_out, r173_out);
	reg32 r174 (rst, clk, r173_out, r174_out);
	reg32 r175 (rst, clk, r174_out, r175_out);
	reg32 r176 (rst, clk, r175_out, r176_out);
	reg32 r177 (rst, clk, r176_out, r177_out);
	reg32 r178 (rst, clk, r177_out, r178_out);
	reg32 r179 (rst, clk, r178_out, r179_out);
	reg32 r180 (rst, clk, r179_out, r180_out);
	reg32 r181 (rst, clk, r180_out, r181_out);
	reg32 r182 (rst, clk, r181_out, r182_out);
	reg32 r183 (rst, clk, r182_out, r183_out);
	reg32 r184 (rst, clk, r183_out, r184_out);
	reg32 r185 (rst, clk, r184_out, r185_out);
	reg32 r186 (rst, clk, r185_out, r186_out);
	reg32 r187 (rst, clk, r186_out, r187_out);
	reg32 r188 (rst, clk, r187_out, r188_out);
	reg32 r189 (rst, clk, r188_out, r189_out);
	reg32 r190 (rst, clk, r189_out, r190_out);
	reg32 r191 (rst, clk, r190_out, r191_out);
	reg32 r192 (rst, clk, r191_out, r192_out);
	reg32 r193 (rst, clk, r192_out, r193_out);
	reg32 r194 (rst, clk, r193_out, r194_out);
	reg32 r195 (rst, clk, r194_out, r195_out);
	reg32 r196 (rst, clk, r195_out, r196_out);
	reg32 r197 (rst, clk, r196_out, r197_out);
	reg32 r198 (rst, clk, r197_out, r198_out);
	reg32 r199 (rst, clk, r198_out, r199_out);
	reg32 r200 (rst, clk, r199_out, r200_out);
	reg32 r201 (rst, clk, r200_out, r201_out);
	reg32 r202 (rst, clk, r201_out, r202_out);
	reg32 r203 (rst, clk, r202_out, r203_out);
	reg32 r204 (rst, clk, r203_out, r204_out);
	reg32 r205 (rst, clk, r204_out, r205_out);
	reg32 r206 (rst, clk, r205_out, r206_out);
	reg32 r207 (rst, clk, r206_out, r207_out);
	reg32 r208 (rst, clk, r207_out, r208_out);
	reg32 r209 (rst, clk, r208_out, r209_out);
	reg32 r210 (rst, clk, r209_out, r210_out);
	reg32 r211 (rst, clk, r210_out, r211_out);
	reg32 r212 (rst, clk, r211_out, r212_out);
	reg32 r213 (rst, clk, r212_out, r213_out);
	reg32 r214 (rst, clk, r213_out, r214_out);
	reg32 r215 (rst, clk, r214_out, r215_out);
	reg32 r216 (rst, clk, r215_out, r216_out);
	reg32 r217 (rst, clk, r216_out, r217_out);
	reg32 r218 (rst, clk, r217_out, r218_out);
	reg32 r219 (rst, clk, r218_out, r219_out);
	reg32 r220 (rst, clk, r219_out, r220_out);
	reg32 r221 (rst, clk, r220_out, r221_out);
	reg32 r222 (rst, clk, r221_out, r222_out);
	reg32 r223 (rst, clk, r222_out, r223_out);
	reg32 r224 (rst, clk, r223_out, r224_out);
	reg32 r225 (rst, clk, r224_out, r225_out);
	reg32 r226 (rst, clk, r225_out, r226_out);
	reg32 r227 (rst, clk, r226_out, r227_out);
	reg32 r228 (rst, clk, r227_out, r228_out);
	reg32 r229 (rst, clk, r228_out, r229_out);
	reg32 r230 (rst, clk, r229_out, r230_out);
	reg32 r231 (rst, clk, r230_out, r231_out);
	reg32 r232 (rst, clk, r231_out, r232_out);
	reg32 r233 (rst, clk, r232_out, r233_out);
	reg32 r234 (rst, clk, r233_out, r234_out);
	reg32 r235 (rst, clk, r234_out, r235_out);
	reg32 r236 (rst, clk, r235_out, r236_out);
	reg32 r237 (rst, clk, r236_out, r237_out);
	reg32 r238 (rst, clk, r237_out, r238_out);
	reg32 r239 (rst, clk, r238_out, r239_out);
	reg32 r240 (rst, clk, r239_out, r240_out);
	reg32 r241 (rst, clk, r240_out, r241_out);
	reg32 r242 (rst, clk, r241_out, r242_out);
	reg32 r243 (rst, clk, r242_out, r243_out);
	reg32 r244 (rst, clk, r243_out, r244_out);
	reg32 r245 (rst, clk, r244_out, r245_out);
	reg32 r246 (rst, clk, r245_out, r246_out);
	reg32 r247 (rst, clk, r246_out, r247_out);
	reg32 r248 (rst, clk, r247_out, r248_out);
	reg32 r249 (rst, clk, r248_out, r249_out);
	reg32 r250 (rst, clk, r249_out, r250_out);
	reg32 r251 (rst, clk, r250_out, r251_out);
	reg32 r252 (rst, clk, r251_out, r252_out);
	reg32 r253 (rst, clk, r252_out, r253_out);
	reg32 r254 (rst, clk, r253_out, r254_out);
	reg32 r255 (rst, clk, r254_out, r255_out);
	reg32 r256 (rst, clk, r255_out, r256_out);
	reg32 r257 (rst, clk, r256_out, r257_out);
	reg32 r258 (rst, clk, r257_out, r258_out);
	reg32 r259 (rst, clk, r258_out, r259_out);
	reg32 r260 (rst, clk, r259_out, r260_out);
	reg32 r261 (rst, clk, r260_out, r261_out);
	reg32 r262 (rst, clk, r261_out, r262_out);
	reg32 r263 (rst, clk, r262_out, r263_out);
	reg32 r264 (rst, clk, r263_out, r264_out);
	reg32 r265 (rst, clk, r264_out, r265_out);
	reg32 r266 (rst, clk, r265_out, r266_out);
	reg32 r267 (rst, clk, r266_out, r267_out);
	reg32 r268 (rst, clk, r267_out, r268_out);
	reg32 r269 (rst, clk, r268_out, r269_out);
	reg32 r270 (rst, clk, r269_out, r270_out);
	reg32 r271 (rst, clk, r270_out, r271_out);
	reg32 r272 (rst, clk, r271_out, r272_out);
	reg32 r273 (rst, clk, r272_out, r273_out);
	reg32 r274 (rst, clk, r273_out, r274_out);
	reg32 r275 (rst, clk, r274_out, r275_out);
	reg32 r276 (rst, clk, r275_out, r276_out);
	reg32 r277 (rst, clk, r276_out, r277_out);
	reg32 r278 (rst, clk, r277_out, r278_out);
	reg32 r279 (rst, clk, r278_out, r279_out);
	reg32 r280 (rst, clk, r279_out, r280_out);
	reg32 r281 (rst, clk, r280_out, r281_out);
	reg32 r282 (rst, clk, r281_out, r282_out);
	reg32 r283 (rst, clk, r282_out, r283_out);
	reg32 r284 (rst, clk, r283_out, r284_out);
	reg32 r285 (rst, clk, r284_out, r285_out);
	reg32 r286 (rst, clk, r285_out, r286_out);
	reg32 r287 (rst, clk, r286_out, r287_out);
	reg32 r288 (rst, clk, r287_out, r288_out);
	reg32 r289 (rst, clk, r288_out, r289_out);
	reg32 r290 (rst, clk, r289_out, r290_out);
	reg32 r291 (rst, clk, r290_out, r291_out);
	reg32 r292 (rst, clk, r291_out, r292_out);
	reg32 r293 (rst, clk, r292_out, r293_out);
	reg32 r294 (rst, clk, r293_out, r294_out);
	reg32 r295 (rst, clk, r294_out, r295_out);
	reg32 r296 (rst, clk, r295_out, r296_out);
	reg32 r297 (rst, clk, r296_out, r297_out);
	reg32 r298 (rst, clk, r297_out, r298_out);
	reg32 r299 (rst, clk, r298_out, r299_out);
	reg32 r300 (rst, clk, r299_out, r300_out);
	reg32 r301 (rst, clk, r300_out, r301_out);
	reg32 r302 (rst, clk, r301_out, r302_out);
	reg32 r303 (rst, clk, r302_out, r303_out);
	reg32 r304 (rst, clk, r303_out, r304_out);
	reg32 r305 (rst, clk, r304_out, r305_out);
	reg32 r306 (rst, clk, r305_out, r306_out);
	reg32 r307 (rst, clk, r306_out, r307_out);
	reg32 r308 (rst, clk, r307_out, r308_out);
	reg32 r309 (rst, clk, r308_out, r309_out);
	reg32 r310 (rst, clk, r309_out, r310_out);
	reg32 r311 (rst, clk, r310_out, r311_out);
	reg32 r312 (rst, clk, r311_out, r312_out);
	reg32 r313 (rst, clk, r312_out, r313_out);
	reg32 r314 (rst, clk, r313_out, r314_out);
	reg32 r315 (rst, clk, r314_out, r315_out);
	reg32 r316 (rst, clk, r315_out, r316_out);
	reg32 r317 (rst, clk, r316_out, r317_out);
	reg32 r318 (rst, clk, r317_out, r318_out);
	reg32 r319 (rst, clk, r318_out, r319_out);
	reg32 r320 (rst, clk, r319_out, r320_out);
	reg32 r321 (rst, clk, r320_out, r321_out);
	reg32 r322 (rst, clk, r321_out, r322_out);
	reg32 r323 (rst, clk, r322_out, r323_out);
	reg32 r324 (rst, clk, r323_out, r324_out);
	reg32 r325 (rst, clk, r324_out, r325_out);
	reg32 r326 (rst, clk, r325_out, r326_out);
	reg32 r327 (rst, clk, r326_out, r327_out);
	reg32 r328 (rst, clk, r327_out, r328_out);
	reg32 r329 (rst, clk, r328_out, r329_out);
	reg32 r330 (rst, clk, r329_out, r330_out);
	reg32 r331 (rst, clk, r330_out, r331_out);
	reg32 r332 (rst, clk, r331_out, r332_out);
	reg32 r333 (rst, clk, r332_out, r333_out);
	reg32 r334 (rst, clk, r333_out, r334_out);
	reg32 r335 (rst, clk, r334_out, r335_out);
	reg32 r336 (rst, clk, r335_out, r336_out);
	reg32 r337 (rst, clk, r336_out, r337_out);
	reg32 r338 (rst, clk, r337_out, r338_out);
	reg32 r339 (rst, clk, r338_out, r339_out);
	reg32 r340 (rst, clk, r339_out, r340_out);
	reg32 r341 (rst, clk, r340_out, r341_out);
	reg32 r342 (rst, clk, r341_out, r342_out);
	reg32 r343 (rst, clk, r342_out, r343_out);
	reg32 r344 (rst, clk, r343_out, r344_out);
	reg32 r345 (rst, clk, r344_out, r345_out);
	reg32 r346 (rst, clk, r345_out, r346_out);
	reg32 r347 (rst, clk, r346_out, r347_out);
	reg32 r348 (rst, clk, r347_out, r348_out);
	reg32 r349 (rst, clk, r348_out, r349_out);
	reg32 r350 (rst, clk, r349_out, r350_out);
	reg32 r351 (rst, clk, r350_out, r351_out);
	reg32 r352 (rst, clk, r351_out, r352_out);
	reg32 r353 (rst, clk, r352_out, r353_out);
	reg32 r354 (rst, clk, r353_out, r354_out);
	reg32 r355 (rst, clk, r354_out, r355_out);
	reg32 r356 (rst, clk, r355_out, r356_out);
	reg32 r357 (rst, clk, r356_out, r357_out);
	reg32 r358 (rst, clk, r357_out, r358_out);
	reg32 r359 (rst, clk, r358_out, r359_out);
	reg32 r360 (rst, clk, r359_out, r360_out);
	reg32 r361 (rst, clk, r360_out, r361_out);
	reg32 r362 (rst, clk, r361_out, r362_out);
	reg32 r363 (rst, clk, r362_out, r363_out);
	reg32 r364 (rst, clk, r363_out, r364_out);
	reg32 r365 (rst, clk, r364_out, r365_out);
	reg32 r366 (rst, clk, r365_out, r366_out);
	reg32 r367 (rst, clk, r366_out, r367_out);
	reg32 r368 (rst, clk, r367_out, r368_out);
	reg32 r369 (rst, clk, r368_out, r369_out);
	reg32 r370 (rst, clk, r369_out, r370_out);
	reg32 r371 (rst, clk, r370_out, r371_out);
	reg32 r372 (rst, clk, r371_out, r372_out);
	reg32 r373 (rst, clk, r372_out, r373_out);
	reg32 r374 (rst, clk, r373_out, r374_out);
	reg32 r375 (rst, clk, r374_out, r375_out);
	reg32 r376 (rst, clk, r375_out, r376_out);
	reg32 r377 (rst, clk, r376_out, r377_out);
	reg32 r378 (rst, clk, r377_out, r378_out);
	reg32 r379 (rst, clk, r378_out, r379_out);
	reg32 r380 (rst, clk, r379_out, r380_out);
	reg32 r381 (rst, clk, r380_out, r381_out);
	reg32 r382 (rst, clk, r381_out, r382_out);
	reg32 r383 (rst, clk, r382_out, r383_out);
	reg32 r384 (rst, clk, r383_out, r384_out);
	reg32 r385 (rst, clk, r384_out, r385_out);
	reg32 r386 (rst, clk, r385_out, r386_out);
	reg32 r387 (rst, clk, r386_out, r387_out);
	reg32 r388 (rst, clk, r387_out, r388_out);
	reg32 r389 (rst, clk, r388_out, r389_out);
	reg32 r390 (rst, clk, r389_out, r390_out);
	reg32 r391 (rst, clk, r390_out, r391_out);
	reg32 r392 (rst, clk, r391_out, r392_out);
	reg32 r393 (rst, clk, r392_out, r393_out);
	reg32 r394 (rst, clk, r393_out, r394_out);
	reg32 r395 (rst, clk, r394_out, r395_out);
	reg32 r396 (rst, clk, r395_out, r396_out);
	reg32 r397 (rst, clk, r396_out, r397_out);
	reg32 r398 (rst, clk, r397_out, r398_out);
	reg32 r399 (rst, clk, r398_out, r399_out);
	reg32 r400 (rst, clk, r399_out, r400_out);
	reg32 r401 (rst, clk, r400_out, r401_out);
	reg32 r402 (rst, clk, r401_out, r402_out);
	reg32 r403 (rst, clk, r402_out, r403_out);
	reg32 r404 (rst, clk, r403_out, r404_out);
	reg32 r405 (rst, clk, r404_out, r405_out);
	reg32 r406 (rst, clk, r405_out, r406_out);
	reg32 r407 (rst, clk, r406_out, r407_out);
	reg32 r408 (rst, clk, r407_out, r408_out);
	reg32 r409 (rst, clk, r408_out, r409_out);
	reg32 r410 (rst, clk, r409_out, r410_out);
	reg32 r411 (rst, clk, r410_out, r411_out);
	reg32 r412 (rst, clk, r411_out, r412_out);
	reg32 r413 (rst, clk, r412_out, r413_out);
	reg32 r414 (rst, clk, r413_out, r414_out);
	reg32 r415 (rst, clk, r414_out, r415_out);
	reg32 r416 (rst, clk, r415_out, r416_out);
	reg32 r417 (rst, clk, r416_out, r417_out);
	reg32 r418 (rst, clk, r417_out, r418_out);
	reg32 r419 (rst, clk, r418_out, r419_out);
	reg32 r420 (rst, clk, r419_out, r420_out);
	reg32 r421 (rst, clk, r420_out, r421_out);
	reg32 r422 (rst, clk, r421_out, r422_out);
	reg32 r423 (rst, clk, r422_out, r423_out);
	reg32 r424 (rst, clk, r423_out, r424_out);
	reg32 r425 (rst, clk, r424_out, r425_out);
	reg32 r426 (rst, clk, r425_out, r426_out);
	reg32 r427 (rst, clk, r426_out, r427_out);
	reg32 r428 (rst, clk, r427_out, r428_out);
	reg32 r429 (rst, clk, r428_out, r429_out);
	reg32 r430 (rst, clk, r429_out, r430_out);
	reg32 r431 (rst, clk, r430_out, r431_out);
	reg32 r432 (rst, clk, r431_out, r432_out);
	reg32 r433 (rst, clk, r432_out, r433_out);
	reg32 r434 (rst, clk, r433_out, r434_out);
	reg32 r435 (rst, clk, r434_out, r435_out);
	reg32 r436 (rst, clk, r435_out, r436_out);
	reg32 r437 (rst, clk, r436_out, r437_out);
	reg32 r438 (rst, clk, r437_out, r438_out);
	reg32 r439 (rst, clk, r438_out, r439_out);
	reg32 r440 (rst, clk, r439_out, r440_out);
	reg32 r441 (rst, clk, r440_out, r441_out);
	reg32 r442 (rst, clk, r441_out, r442_out);
	reg32 r443 (rst, clk, r442_out, r443_out);
	reg32 r444 (rst, clk, r443_out, r444_out);
	reg32 r445 (rst, clk, r444_out, r445_out);
	reg32 r446 (rst, clk, r445_out, r446_out);
	reg32 r447 (rst, clk, r446_out, r447_out);
	reg32 r448 (rst, clk, r447_out, r448_out);
	reg32 r449 (rst, clk, r448_out, r449_out);
	reg32 r450 (rst, clk, r449_out, r450_out);
	reg32 r451 (rst, clk, r450_out, r451_out);
	reg32 r452 (rst, clk, r451_out, r452_out);
	reg32 r453 (rst, clk, r452_out, r453_out);
	reg32 r454 (rst, clk, r453_out, r454_out);
	reg32 r455 (rst, clk, r454_out, r455_out);
	reg32 r456 (rst, clk, r455_out, r456_out);
	reg32 r457 (rst, clk, r456_out, r457_out);
	reg32 r458 (rst, clk, r457_out, r458_out);
	reg32 r459 (rst, clk, r458_out, r459_out);
	reg32 r460 (rst, clk, r459_out, r460_out);
	reg32 r461 (rst, clk, r460_out, r461_out);
	reg32 r462 (rst, clk, r461_out, r462_out);
	reg32 r463 (rst, clk, r462_out, r463_out);
	reg32 r464 (rst, clk, r463_out, r464_out);
	reg32 r465 (rst, clk, r464_out, r465_out);
	reg32 r466 (rst, clk, r465_out, r466_out);
	reg32 r467 (rst, clk, r466_out, r467_out);
	reg32 r468 (rst, clk, r467_out, r468_out);
	reg32 r469 (rst, clk, r468_out, r469_out);
	reg32 r470 (rst, clk, r469_out, r470_out);
	reg32 r471 (rst, clk, r470_out, r471_out);
	reg32 r472 (rst, clk, r471_out, r472_out);
	reg32 r473 (rst, clk, r472_out, r473_out);
	reg32 r474 (rst, clk, r473_out, r474_out);
	reg32 r475 (rst, clk, r474_out, r475_out);
	reg32 r476 (rst, clk, r475_out, r476_out);
	reg32 r477 (rst, clk, r476_out, r477_out);
	reg32 r478 (rst, clk, r477_out, r478_out);
	reg32 r479 (rst, clk, r478_out, r479_out);
	reg32 r480 (rst, clk, r479_out, r480_out);
	reg32 r481 (rst, clk, r480_out, r481_out);
	reg32 r482 (rst, clk, r481_out, r482_out);
	reg32 r483 (rst, clk, r482_out, r483_out);
	reg32 r484 (rst, clk, r483_out, r484_out);
	reg32 r485 (rst, clk, r484_out, r485_out);
	reg32 r486 (rst, clk, r485_out, r486_out);
	reg32 r487 (rst, clk, r486_out, r487_out);
	reg32 r488 (rst, clk, r487_out, r488_out);
	reg32 r489 (rst, clk, r488_out, r489_out);
	reg32 r490 (rst, clk, r489_out, r490_out);
	reg32 r491 (rst, clk, r490_out, r491_out);
	reg32 r492 (rst, clk, r491_out, r492_out);
	reg32 r493 (rst, clk, r492_out, r493_out);
	reg32 r494 (rst, clk, r493_out, r494_out);
	reg32 r495 (rst, clk, r494_out, r495_out);
	reg32 r496 (rst, clk, r495_out, r496_out);
	reg32 r497 (rst, clk, r496_out, r497_out);
	reg32 r498 (rst, clk, r497_out, r498_out);
	reg32 r499 (rst, clk, r498_out, r499_out);
	reg32 r500 (rst, clk, r499_out, r500_out);
	reg32 r501 (rst, clk, r500_out, r501_out);
	reg32 r502 (rst, clk, r501_out, r502_out);
	reg32 r503 (rst, clk, r502_out, r503_out);
	reg32 r504 (rst, clk, r503_out, r504_out);
	reg32 r505 (rst, clk, r504_out, r505_out);
	reg32 r506 (rst, clk, r505_out, r506_out);
	reg32 r507 (rst, clk, r506_out, r507_out);
	reg32 r508 (rst, clk, r507_out, r508_out);
	reg32 r509 (rst, clk, r508_out, r509_out);
	reg32 r510 (rst, clk, r509_out, r510_out);
	reg32 r511 (rst, clk, r510_out, r511_out);
	reg32 r512 (rst, clk, r511_out, r512_out);
	reg32 r513 (rst, clk, r512_out, r513_out);
	reg32 r514 (rst, clk, r513_out, r514_out);
	reg32 r515 (rst, clk, r514_out, r515_out);
	reg32 r516 (rst, clk, r515_out, r516_out);
	reg32 r517 (rst, clk, r516_out, r517_out);
	reg32 r518 (rst, clk, r517_out, r518_out);
	reg32 r519 (rst, clk, r518_out, r519_out);
	reg32 r520 (rst, clk, r519_out, r520_out);
	reg32 r521 (rst, clk, r520_out, r521_out);
	reg32 r522 (rst, clk, r521_out, r522_out);
	reg32 r523 (rst, clk, r522_out, r523_out);
	reg32 r524 (rst, clk, r523_out, r524_out);
	reg32 r525 (rst, clk, r524_out, r525_out);
	reg32 r526 (rst, clk, r525_out, r526_out);
	reg32 r527 (rst, clk, r526_out, r527_out);
	reg32 r528 (rst, clk, r527_out, r528_out);
	reg32 r529 (rst, clk, r528_out, r529_out);
	reg32 r530 (rst, clk, r529_out, r530_out);
	reg32 r531 (rst, clk, r530_out, r531_out);
	reg32 r532 (rst, clk, r531_out, r532_out);
	reg32 r533 (rst, clk, r532_out, r533_out);
	reg32 r534 (rst, clk, r533_out, r534_out);
	reg32 r535 (rst, clk, r534_out, r535_out);
	reg32 r536 (rst, clk, r535_out, r536_out);
	reg32 r537 (rst, clk, r536_out, r537_out);
	reg32 r538 (rst, clk, r537_out, r538_out);
	reg32 r539 (rst, clk, r538_out, r539_out);
	reg32 r540 (rst, clk, r539_out, r540_out);
	reg32 r541 (rst, clk, r540_out, r541_out);
	reg32 r542 (rst, clk, r541_out, r542_out);
	reg32 r543 (rst, clk, r542_out, r543_out);
	reg32 r544 (rst, clk, r543_out, r544_out);
	reg32 r545 (rst, clk, r544_out, r545_out);
	reg32 r546 (rst, clk, r545_out, r546_out);
	reg32 r547 (rst, clk, r546_out, r547_out);
	reg32 r548 (rst, clk, r547_out, r548_out);
	reg32 r549 (rst, clk, r548_out, r549_out);
	reg32 r550 (rst, clk, r549_out, r550_out);
	reg32 r551 (rst, clk, r550_out, r551_out);
	reg32 r552 (rst, clk, r551_out, r552_out);
	reg32 r553 (rst, clk, r552_out, r553_out);
	reg32 r554 (rst, clk, r553_out, r554_out);
	reg32 r555 (rst, clk, r554_out, r555_out);
	reg32 r556 (rst, clk, r555_out, r556_out);
	reg32 r557 (rst, clk, r556_out, r557_out);
	reg32 r558 (rst, clk, r557_out, r558_out);
	reg32 r559 (rst, clk, r558_out, r559_out);
	reg32 r560 (rst, clk, r559_out, r560_out);
	reg32 r561 (rst, clk, r560_out, r561_out);
	reg32 r562 (rst, clk, r561_out, r562_out);
	reg32 r563 (rst, clk, r562_out, r563_out);
	reg32 r564 (rst, clk, r563_out, r564_out);
	reg32 r565 (rst, clk, r564_out, r565_out);
	reg32 r566 (rst, clk, r565_out, r566_out);
	reg32 r567 (rst, clk, r566_out, r567_out);
	reg32 r568 (rst, clk, r567_out, r568_out);
	reg32 r569 (rst, clk, r568_out, r569_out);
	reg32 r570 (rst, clk, r569_out, r570_out);
	reg32 r571 (rst, clk, r570_out, r571_out);
	reg32 r572 (rst, clk, r571_out, r572_out);
	reg32 r573 (rst, clk, r572_out, r573_out);
	reg32 r574 (rst, clk, r573_out, r574_out);
	reg32 r575 (rst, clk, r574_out, r575_out);
	reg32 r576 (rst, clk, r575_out, r576_out);
	reg32 r577 (rst, clk, r576_out, r577_out);
	reg32 r578 (rst, clk, r577_out, r578_out);
	reg32 r579 (rst, clk, r578_out, r579_out);
	reg32 r580 (rst, clk, r579_out, r580_out);
	reg32 r581 (rst, clk, r580_out, r581_out);
	reg32 r582 (rst, clk, r581_out, r582_out);
	reg32 r583 (rst, clk, r582_out, r583_out);
	reg32 r584 (rst, clk, r583_out, r584_out);
	reg32 r585 (rst, clk, r584_out, r585_out);
	reg32 r586 (rst, clk, r585_out, r586_out);
	reg32 r587 (rst, clk, r586_out, r587_out);
	reg32 r588 (rst, clk, r587_out, r588_out);
	reg32 r589 (rst, clk, r588_out, r589_out);
	reg32 r590 (rst, clk, r589_out, r590_out);
	reg32 r591 (rst, clk, r590_out, r591_out);
	reg32 r592 (rst, clk, r591_out, r592_out);
	reg32 r593 (rst, clk, r592_out, r593_out);
	reg32 r594 (rst, clk, r593_out, r594_out);
	reg32 r595 (rst, clk, r594_out, r595_out);
	reg32 r596 (rst, clk, r595_out, r596_out);
	reg32 r597 (rst, clk, r596_out, r597_out);
	reg32 r598 (rst, clk, r597_out, r598_out);
	reg32 r599 (rst, clk, r598_out, r599_out);
	reg32 r600 (rst, clk, r599_out, r600_out);
	reg32 r601 (rst, clk, r600_out, r601_out);
	reg32 r602 (rst, clk, r601_out, r602_out);
	reg32 r603 (rst, clk, r602_out, r603_out);
	reg32 r604 (rst, clk, r603_out, r604_out);
	reg32 r605 (rst, clk, r604_out, r605_out);
	reg32 r606 (rst, clk, r605_out, r606_out);
	reg32 r607 (rst, clk, r606_out, r607_out);
	reg32 r608 (rst, clk, r607_out, r608_out);
	reg32 r609 (rst, clk, r608_out, r609_out);
	reg32 r610 (rst, clk, r609_out, r610_out);
	reg32 r611 (rst, clk, r610_out, r611_out);
	reg32 r612 (rst, clk, r611_out, r612_out);
	reg32 r613 (rst, clk, r612_out, r613_out);
	reg32 r614 (rst, clk, r613_out, r614_out);
	reg32 r615 (rst, clk, r614_out, r615_out);
	reg32 r616 (rst, clk, r615_out, r616_out);
	reg32 r617 (rst, clk, r616_out, r617_out);
	reg32 r618 (rst, clk, r617_out, r618_out);
	reg32 r619 (rst, clk, r618_out, r619_out);
	reg32 r620 (rst, clk, r619_out, r620_out);
	reg32 r621 (rst, clk, r620_out, r621_out);
	reg32 r622 (rst, clk, r621_out, r622_out);
	reg32 r623 (rst, clk, r622_out, r623_out);
	reg32 r624 (rst, clk, r623_out, r624_out);
	reg32 r625 (rst, clk, r624_out, r625_out);
	reg32 r626 (rst, clk, r625_out, r626_out);
	reg32 r627 (rst, clk, r626_out, r627_out);
	reg32 r628 (rst, clk, r627_out, r628_out);
	reg32 r629 (rst, clk, r628_out, r629_out);
	reg32 r630 (rst, clk, r629_out, r630_out);
	reg32 r631 (rst, clk, r630_out, r631_out);
	reg32 r632 (rst, clk, r631_out, r632_out);
	reg32 r633 (rst, clk, r632_out, r633_out);
	reg32 r634 (rst, clk, r633_out, r634_out);
	reg32 r635 (rst, clk, r634_out, r635_out);
	reg32 r636 (rst, clk, r635_out, r636_out);
	reg32 r637 (rst, clk, r636_out, r637_out);
	reg32 r638 (rst, clk, r637_out, r638_out);
	reg32 r639 (rst, clk, r638_out, r639_out);
	reg32 r640 (rst, clk, r639_out, r640_out);
	reg32 r641 (rst, clk, r640_out, r641_out);
	reg32 r642 (rst, clk, r641_out, r642_out);
	reg32 r643 (rst, clk, r642_out, r643_out);
	reg32 r644 (rst, clk, r643_out, r644_out);
	reg32 r645 (rst, clk, r644_out, r645_out);
	reg32 r646 (rst, clk, r645_out, r646_out);
	reg32 r647 (rst, clk, r646_out, r647_out);
	reg32 r648 (rst, clk, r647_out, r648_out);
	reg32 r649 (rst, clk, r648_out, r649_out);
	reg32 r650 (rst, clk, r649_out, r650_out);
	reg32 r651 (rst, clk, r650_out, r651_out);
	reg32 r652 (rst, clk, r651_out, r652_out);
	reg32 r653 (rst, clk, r652_out, r653_out);
	reg32 r654 (rst, clk, r653_out, r654_out);
	reg32 r655 (rst, clk, r654_out, r655_out);
	reg32 r656 (rst, clk, r655_out, r656_out);
	reg32 r657 (rst, clk, r656_out, r657_out);
	reg32 r658 (rst, clk, r657_out, r658_out);
	reg32 r659 (rst, clk, r658_out, r659_out);
	reg32 r660 (rst, clk, r659_out, r660_out);
	reg32 r661 (rst, clk, r660_out, r661_out);
	reg32 r662 (rst, clk, r661_out, r662_out);
	reg32 r663 (rst, clk, r662_out, r663_out);
	reg32 r664 (rst, clk, r663_out, r664_out);
	reg32 r665 (rst, clk, r664_out, r665_out);
	reg32 r666 (rst, clk, r665_out, r666_out);
	reg32 r667 (rst, clk, r666_out, r667_out);
	reg32 r668 (rst, clk, r667_out, r668_out);
	reg32 r669 (rst, clk, r668_out, r669_out);
	reg32 r670 (rst, clk, r669_out, r670_out);
	reg32 r671 (rst, clk, r670_out, r671_out);
	reg32 r672 (rst, clk, r671_out, r672_out);
	reg32 r673 (rst, clk, r672_out, r673_out);
	reg32 r674 (rst, clk, r673_out, r674_out);
	reg32 r675 (rst, clk, r674_out, r675_out);
	reg32 r676 (rst, clk, r675_out, r676_out);
	reg32 r677 (rst, clk, r676_out, r677_out);
	reg32 r678 (rst, clk, r677_out, r678_out);
	reg32 r679 (rst, clk, r678_out, r679_out);
	reg32 r680 (rst, clk, r679_out, r680_out);
	reg32 r681 (rst, clk, r680_out, r681_out);
	reg32 r682 (rst, clk, r681_out, r682_out);
	reg32 r683 (rst, clk, r682_out, r683_out);
	reg32 r684 (rst, clk, r683_out, r684_out);
	reg32 r685 (rst, clk, r684_out, r685_out);
	reg32 r686 (rst, clk, r685_out, r686_out);
	reg32 r687 (rst, clk, r686_out, r687_out);
	reg32 r688 (rst, clk, r687_out, r688_out);
	reg32 r689 (rst, clk, r688_out, r689_out);
	reg32 r690 (rst, clk, r689_out, r690_out);
	reg32 r691 (rst, clk, r690_out, r691_out);
	reg32 r692 (rst, clk, r691_out, r692_out);
	reg32 r693 (rst, clk, r692_out, r693_out);
	reg32 r694 (rst, clk, r693_out, r694_out);
	reg32 r695 (rst, clk, r694_out, r695_out);
	reg32 r696 (rst, clk, r695_out, r696_out);
	reg32 r697 (rst, clk, r696_out, r697_out);
	reg32 r698 (rst, clk, r697_out, r698_out);
	reg32 r699 (rst, clk, r698_out, r699_out);
	reg32 r700 (rst, clk, r699_out, r700_out);
	reg32 r701 (rst, clk, r700_out, r701_out);
	reg32 r702 (rst, clk, r701_out, r702_out);
	reg32 r703 (rst, clk, r702_out, r703_out);
	reg32 r704 (rst, clk, r703_out, r704_out);
	reg32 r705 (rst, clk, r704_out, r705_out);
	reg32 r706 (rst, clk, r705_out, r706_out);
	reg32 r707 (rst, clk, r706_out, r707_out);
	reg32 r708 (rst, clk, r707_out, r708_out);
	reg32 r709 (rst, clk, r708_out, r709_out);
	reg32 r710 (rst, clk, r709_out, r710_out);
	reg32 r711 (rst, clk, r710_out, r711_out);
	reg32 r712 (rst, clk, r711_out, r712_out);
	reg32 r713 (rst, clk, r712_out, r713_out);
	reg32 r714 (rst, clk, r713_out, r714_out);
	reg32 r715 (rst, clk, r714_out, r715_out);
	reg32 r716 (rst, clk, r715_out, r716_out);
	reg32 r717 (rst, clk, r716_out, r717_out);
	reg32 r718 (rst, clk, r717_out, r718_out);
	reg32 r719 (rst, clk, r718_out, r719_out);
	reg32 r720 (rst, clk, r719_out, r720_out);
	reg32 r721 (rst, clk, r720_out, r721_out);
	reg32 r722 (rst, clk, r721_out, r722_out);
	reg32 r723 (rst, clk, r722_out, r723_out);
	reg32 r724 (rst, clk, r723_out, r724_out);
	reg32 r725 (rst, clk, r724_out, r725_out);
	reg32 r726 (rst, clk, r725_out, r726_out);
	reg32 r727 (rst, clk, r726_out, r727_out);
	reg32 r728 (rst, clk, r727_out, r728_out);
	reg32 r729 (rst, clk, r728_out, r729_out);
	reg32 r730 (rst, clk, r729_out, r730_out);
	reg32 r731 (rst, clk, r730_out, r731_out);
	reg32 r732 (rst, clk, r731_out, r732_out);
	reg32 r733 (rst, clk, r732_out, r733_out);
	reg32 r734 (rst, clk, r733_out, r734_out);
	reg32 r735 (rst, clk, r734_out, r735_out);
	reg32 r736 (rst, clk, r735_out, r736_out);
	reg32 r737 (rst, clk, r736_out, r737_out);
	reg32 r738 (rst, clk, r737_out, r738_out);
	reg32 r739 (rst, clk, r738_out, r739_out);
	reg32 r740 (rst, clk, r739_out, r740_out);
	reg32 r741 (rst, clk, r740_out, r741_out);
	reg32 r742 (rst, clk, r741_out, r742_out);
	reg32 r743 (rst, clk, r742_out, r743_out);
	reg32 r744 (rst, clk, r743_out, r744_out);
	reg32 r745 (rst, clk, r744_out, r745_out);
	reg32 r746 (rst, clk, r745_out, r746_out);
	reg32 r747 (rst, clk, r746_out, r747_out);
	reg32 r748 (rst, clk, r747_out, r748_out);
	reg32 r749 (rst, clk, r748_out, r749_out);
	reg32 r750 (rst, clk, r749_out, r750_out);
	reg32 r751 (rst, clk, r750_out, r751_out);
	reg32 r752 (rst, clk, r751_out, r752_out);
	reg32 r753 (rst, clk, r752_out, r753_out);
	reg32 r754 (rst, clk, r753_out, r754_out);
	reg32 r755 (rst, clk, r754_out, r755_out);
	reg32 r756 (rst, clk, r755_out, r756_out);
	reg32 r757 (rst, clk, r756_out, r757_out);
	reg32 r758 (rst, clk, r757_out, r758_out);
	reg32 r759 (rst, clk, r758_out, r759_out);
	reg32 r760 (rst, clk, r759_out, r760_out);
	reg32 r761 (rst, clk, r760_out, r761_out);
	reg32 r762 (rst, clk, r761_out, r762_out);
	reg32 r763 (rst, clk, r762_out, r763_out);
	reg32 r764 (rst, clk, r763_out, r764_out);
	reg32 r765 (rst, clk, r764_out, r765_out);
	reg32 r766 (rst, clk, r765_out, r766_out);
	reg32 r767 (rst, clk, r766_out, r767_out);
	reg32 r768 (rst, clk, r767_out, r768_out);
	reg32 r769 (rst, clk, r768_out, r769_out);
	reg32 r770 (rst, clk, r769_out, r770_out);
	reg32 r771 (rst, clk, r770_out, r771_out);
	reg32 r772 (rst, clk, r771_out, r772_out);
	reg32 r773 (rst, clk, r772_out, r773_out);
	reg32 r774 (rst, clk, r773_out, r774_out);
	reg32 r775 (rst, clk, r774_out, r775_out);
	reg32 r776 (rst, clk, r775_out, r776_out);
	reg32 r777 (rst, clk, r776_out, r777_out);
	reg32 r778 (rst, clk, r777_out, r778_out);
	reg32 r779 (rst, clk, r778_out, r779_out);
	reg32 r780 (rst, clk, r779_out, r780_out);
	reg32 r781 (rst, clk, r780_out, r781_out);
	reg32 r782 (rst, clk, r781_out, r782_out);
	reg32 r783 (rst, clk, r782_out, r783_out);
	reg32 r784 (rst, clk, r783_out, r784_out);
	reg32 r785 (rst, clk, r784_out, r785_out);
	reg32 r786 (rst, clk, r785_out, r786_out);
	reg32 r787 (rst, clk, r786_out, r787_out);
	reg32 r788 (rst, clk, r787_out, r788_out);
	reg32 r789 (rst, clk, r788_out, r789_out);
	reg32 r790 (rst, clk, r789_out, r790_out);
	reg32 r791 (rst, clk, r790_out, r791_out);
	reg32 r792 (rst, clk, r791_out, r792_out);
	reg32 r793 (rst, clk, r792_out, r793_out);
	reg32 r794 (rst, clk, r793_out, r794_out);
	reg32 r795 (rst, clk, r794_out, r795_out);
	reg32 r796 (rst, clk, r795_out, r796_out);
	reg32 r797 (rst, clk, r796_out, r797_out);
	reg32 r798 (rst, clk, r797_out, r798_out);
	reg32 r799 (rst, clk, r798_out, r799_out);
	reg32 r800 (rst, clk, r799_out, r800_out);
	reg32 r801 (rst, clk, r800_out, r801_out);
	reg32 r802 (rst, clk, r801_out, r802_out);
	reg32 r803 (rst, clk, r802_out, r803_out);
	reg32 r804 (rst, clk, r803_out, r804_out);
	reg32 r805 (rst, clk, r804_out, r805_out);
	reg32 r806 (rst, clk, r805_out, r806_out);
	reg32 r807 (rst, clk, r806_out, r807_out);
	reg32 r808 (rst, clk, r807_out, r808_out);
	reg32 r809 (rst, clk, r808_out, r809_out);
	reg32 r810 (rst, clk, r809_out, r810_out);
	reg32 r811 (rst, clk, r810_out, r811_out);
	reg32 r812 (rst, clk, r811_out, r812_out);
	reg32 r813 (rst, clk, r812_out, r813_out);
	reg32 r814 (rst, clk, r813_out, r814_out);
	reg32 r815 (rst, clk, r814_out, r815_out);
	reg32 r816 (rst, clk, r815_out, r816_out);
	reg32 r817 (rst, clk, r816_out, r817_out);
	reg32 r818 (rst, clk, r817_out, r818_out);
	reg32 r819 (rst, clk, r818_out, r819_out);
	reg32 r820 (rst, clk, r819_out, r820_out);
	reg32 r821 (rst, clk, r820_out, r821_out);
	reg32 r822 (rst, clk, r821_out, r822_out);
	reg32 r823 (rst, clk, r822_out, r823_out);
	reg32 r824 (rst, clk, r823_out, r824_out);
	reg32 r825 (rst, clk, r824_out, r825_out);
	reg32 r826 (rst, clk, r825_out, r826_out);
	reg32 r827 (rst, clk, r826_out, r827_out);
	reg32 r828 (rst, clk, r827_out, r828_out);
	reg32 r829 (rst, clk, r828_out, r829_out);
	reg32 r830 (rst, clk, r829_out, r830_out);
	reg32 r831 (rst, clk, r830_out, r831_out);
	reg32 r832 (rst, clk, r831_out, r832_out);
	reg32 r833 (rst, clk, r832_out, r833_out);
	reg32 r834 (rst, clk, r833_out, r834_out);
	reg32 r835 (rst, clk, r834_out, r835_out);
	reg32 r836 (rst, clk, r835_out, r836_out);
	reg32 r837 (rst, clk, r836_out, r837_out);
	reg32 r838 (rst, clk, r837_out, r838_out);
	reg32 r839 (rst, clk, r838_out, r839_out);
	reg32 r840 (rst, clk, r839_out, r840_out);
	reg32 r841 (rst, clk, r840_out, r841_out);
	reg32 r842 (rst, clk, r841_out, r842_out);
	reg32 r843 (rst, clk, r842_out, r843_out);
	reg32 r844 (rst, clk, r843_out, r844_out);
	reg32 r845 (rst, clk, r844_out, r845_out);
	reg32 r846 (rst, clk, r845_out, r846_out);
	reg32 r847 (rst, clk, r846_out, r847_out);
	reg32 r848 (rst, clk, r847_out, r848_out);
	reg32 r849 (rst, clk, r848_out, r849_out);
	reg32 r850 (rst, clk, r849_out, r850_out);
	reg32 r851 (rst, clk, r850_out, r851_out);
	reg32 r852 (rst, clk, r851_out, r852_out);
	reg32 r853 (rst, clk, r852_out, r853_out);
	reg32 r854 (rst, clk, r853_out, r854_out);
	reg32 r855 (rst, clk, r854_out, r855_out);
	reg32 r856 (rst, clk, r855_out, r856_out);
	reg32 r857 (rst, clk, r856_out, r857_out);
	reg32 r858 (rst, clk, r857_out, r858_out);
	reg32 r859 (rst, clk, r858_out, r859_out);
	reg32 r860 (rst, clk, r859_out, r860_out);
	reg32 r861 (rst, clk, r860_out, r861_out);
	reg32 r862 (rst, clk, r861_out, r862_out);
	reg32 r863 (rst, clk, r862_out, r863_out);
	reg32 r864 (rst, clk, r863_out, r864_out);
	reg32 r865 (rst, clk, r864_out, r865_out);
	reg32 r866 (rst, clk, r865_out, r866_out);
	reg32 r867 (rst, clk, r866_out, r867_out);
	reg32 r868 (rst, clk, r867_out, r868_out);
	reg32 r869 (rst, clk, r868_out, r869_out);
	reg32 r870 (rst, clk, r869_out, r870_out);
	reg32 r871 (rst, clk, r870_out, r871_out);
	reg32 r872 (rst, clk, r871_out, r872_out);
	reg32 r873 (rst, clk, r872_out, r873_out);
	reg32 r874 (rst, clk, r873_out, r874_out);
	reg32 r875 (rst, clk, r874_out, r875_out);
	reg32 r876 (rst, clk, r875_out, r876_out);
	reg32 r877 (rst, clk, r876_out, r877_out);
	reg32 r878 (rst, clk, r877_out, r878_out);
	reg32 r879 (rst, clk, r878_out, r879_out);
	reg32 r880 (rst, clk, r879_out, r880_out);
	reg32 r881 (rst, clk, r880_out, r881_out);
	reg32 r882 (rst, clk, r881_out, r882_out);
	reg32 r883 (rst, clk, r882_out, r883_out);
	reg32 r884 (rst, clk, r883_out, r884_out);
	reg32 r885 (rst, clk, r884_out, r885_out);
	reg32 r886 (rst, clk, r885_out, r886_out);
	reg32 r887 (rst, clk, r886_out, r887_out);
	reg32 r888 (rst, clk, r887_out, r888_out);
	reg32 r889 (rst, clk, r888_out, r889_out);
	reg32 r890 (rst, clk, r889_out, r890_out);
	reg32 r891 (rst, clk, r890_out, r891_out);
	reg32 r892 (rst, clk, r891_out, r892_out);
	reg32 r893 (rst, clk, r892_out, r893_out);
	reg32 r894 (rst, clk, r893_out, r894_out);
	reg32 r895 (rst, clk, r894_out, r895_out);
	reg32 r896 (rst, clk, r895_out, r896_out);
	reg32 r897 (rst, clk, r896_out, r897_out);
	reg32 r898 (rst, clk, r897_out, r898_out);
	reg32 r899 (rst, clk, r898_out, r899_out);
	reg32 r900 (rst, clk, r899_out, r900_out);
	reg32 r901 (rst, clk, r900_out, r901_out);
	reg32 r902 (rst, clk, r901_out, r902_out);
	reg32 r903 (rst, clk, r902_out, r903_out);
	reg32 r904 (rst, clk, r903_out, r904_out);
	reg32 r905 (rst, clk, r904_out, r905_out);
	reg32 r906 (rst, clk, r905_out, r906_out);
	reg32 r907 (rst, clk, r906_out, r907_out);
	reg32 r908 (rst, clk, r907_out, r908_out);
	reg32 r909 (rst, clk, r908_out, r909_out);
	reg32 r910 (rst, clk, r909_out, r910_out);
	reg32 r911 (rst, clk, r910_out, r911_out);
	reg32 r912 (rst, clk, r911_out, r912_out);
	reg32 r913 (rst, clk, r912_out, r913_out);
	reg32 r914 (rst, clk, r913_out, r914_out);
	reg32 r915 (rst, clk, r914_out, r915_out);
	reg32 r916 (rst, clk, r915_out, r916_out);
	reg32 r917 (rst, clk, r916_out, r917_out);
	reg32 r918 (rst, clk, r917_out, r918_out);
	reg32 r919 (rst, clk, r918_out, r919_out);
	reg32 r920 (rst, clk, r919_out, r920_out);
	reg32 r921 (rst, clk, r920_out, r921_out);
	reg32 r922 (rst, clk, r921_out, r922_out);
	reg32 r923 (rst, clk, r922_out, r923_out);
	reg32 r924 (rst, clk, r923_out, r924_out);
	reg32 r925 (rst, clk, r924_out, r925_out);
	reg32 r926 (rst, clk, r925_out, r926_out);
	reg32 r927 (rst, clk, r926_out, r927_out);
	reg32 r928 (rst, clk, r927_out, r928_out);
	reg32 r929 (rst, clk, r928_out, r929_out);
	reg32 r930 (rst, clk, r929_out, r930_out);
	reg32 r931 (rst, clk, r930_out, r931_out);
	reg32 r932 (rst, clk, r931_out, r932_out);
	reg32 r933 (rst, clk, r932_out, r933_out);
	reg32 r934 (rst, clk, r933_out, r934_out);
	reg32 r935 (rst, clk, r934_out, r935_out);
	reg32 r936 (rst, clk, r935_out, r936_out);
	reg32 r937 (rst, clk, r936_out, r937_out);
	reg32 r938 (rst, clk, r937_out, r938_out);
	reg32 r939 (rst, clk, r938_out, r939_out);
	reg32 r940 (rst, clk, r939_out, r940_out);
	reg32 r941 (rst, clk, r940_out, r941_out);
	reg32 r942 (rst, clk, r941_out, r942_out);
	reg32 r943 (rst, clk, r942_out, r943_out);
	reg32 r944 (rst, clk, r943_out, r944_out);
	reg32 r945 (rst, clk, r944_out, r945_out);
	reg32 r946 (rst, clk, r945_out, r946_out);
	reg32 r947 (rst, clk, r946_out, r947_out);
	reg32 r948 (rst, clk, r947_out, r948_out);
	reg32 r949 (rst, clk, r948_out, r949_out);
	reg32 r950 (rst, clk, r949_out, r950_out);
	reg32 r951 (rst, clk, r950_out, r951_out);
	reg32 r952 (rst, clk, r951_out, r952_out);
	reg32 r953 (rst, clk, r952_out, r953_out);
	reg32 r954 (rst, clk, r953_out, r954_out);
	reg32 r955 (rst, clk, r954_out, r955_out);
	reg32 r956 (rst, clk, r955_out, r956_out);
	reg32 r957 (rst, clk, r956_out, r957_out);
	reg32 r958 (rst, clk, r957_out, r958_out);
	reg32 r959 (rst, clk, r958_out, r959_out);
	reg32 r960 (rst, clk, r959_out, r960_out);
	reg32 r961 (rst, clk, r960_out, r961_out);
	reg32 r962 (rst, clk, r961_out, r962_out);
	reg32 r963 (rst, clk, r962_out, r963_out);
	reg32 r964 (rst, clk, r963_out, r964_out);
	reg32 r965 (rst, clk, r964_out, r965_out);
	reg32 r966 (rst, clk, r965_out, r966_out);
	reg32 r967 (rst, clk, r966_out, r967_out);
	reg32 r968 (rst, clk, r967_out, r968_out);
	reg32 r969 (rst, clk, r968_out, r969_out);
	reg32 r970 (rst, clk, r969_out, r970_out);
	reg32 r971 (rst, clk, r970_out, r971_out);
	reg32 r972 (rst, clk, r971_out, r972_out);
	reg32 r973 (rst, clk, r972_out, r973_out);
	reg32 r974 (rst, clk, r973_out, r974_out);
	reg32 r975 (rst, clk, r974_out, r975_out);
	reg32 r976 (rst, clk, r975_out, r976_out);
	reg32 r977 (rst, clk, r976_out, r977_out);
	reg32 r978 (rst, clk, r977_out, r978_out);
	reg32 r979 (rst, clk, r978_out, r979_out);
	reg32 r980 (rst, clk, r979_out, r980_out);
	reg32 r981 (rst, clk, r980_out, r981_out);
	reg32 r982 (rst, clk, r981_out, r982_out);
	reg32 r983 (rst, clk, r982_out, r983_out);
	reg32 r984 (rst, clk, r983_out, r984_out);
	reg32 r985 (rst, clk, r984_out, r985_out);
	reg32 r986 (rst, clk, r985_out, r986_out);
	reg32 r987 (rst, clk, r986_out, r987_out);
	reg32 r988 (rst, clk, r987_out, r988_out);
	reg32 r989 (rst, clk, r988_out, r989_out);
	reg32 r990 (rst, clk, r989_out, r990_out);
	reg32 r991 (rst, clk, r990_out, r991_out);
	reg32 r992 (rst, clk, r991_out, r992_out);
	reg32 r993 (rst, clk, r992_out, r993_out);
	reg32 r994 (rst, clk, r993_out, r994_out);
	reg32 r995 (rst, clk, r994_out, r995_out);
	reg32 r996 (rst, clk, r995_out, r996_out);
	reg32 r997 (rst, clk, r996_out, r997_out);
	reg32 r998 (rst, clk, r997_out, r998_out);
	reg32 r999 (rst, clk, r998_out, r999_out);
	reg32 r1000 (rst, clk, r999_out, r1000_out);
	reg32 r1001 (rst, clk, r1000_out, r1001_out);
	reg32 r1002 (rst, clk, r1001_out, r1002_out);
	reg32 r1003 (rst, clk, r1002_out, r1003_out);
	reg32 r1004 (rst, clk, r1003_out, r1004_out);
	reg32 r1005 (rst, clk, r1004_out, r1005_out);
	reg32 r1006 (rst, clk, r1005_out, r1006_out);
	reg32 r1007 (rst, clk, r1006_out, r1007_out);
	reg32 r1008 (rst, clk, r1007_out, r1008_out);
	reg32 r1009 (rst, clk, r1008_out, r1009_out);
	reg32 r1010 (rst, clk, r1009_out, r1010_out);
	reg32 r1011 (rst, clk, r1010_out, r1011_out);
	reg32 r1012 (rst, clk, r1011_out, r1012_out);
	reg32 r1013 (rst, clk, r1012_out, r1013_out);
	reg32 r1014 (rst, clk, r1013_out, r1014_out);
	reg32 r1015 (rst, clk, r1014_out, r1015_out);
	reg32 r1016 (rst, clk, r1015_out, r1016_out);
	reg32 r1017 (rst, clk, r1016_out, r1017_out);
	reg32 r1018 (rst, clk, r1017_out, r1018_out);
	reg32 r1019 (rst, clk, r1018_out, r1019_out);
	reg32 r1020 (rst, clk, r1019_out, r1020_out);
	reg32 r1021 (rst, clk, r1020_out, r1021_out);
	reg32 r1022 (rst, clk, r1021_out, r1022_out);
	reg32 r1023 (rst, clk, r1022_out, r1023_out);
	reg32 r1024 (rst, clk, r1023_out, r1024_out);
	reg32 r1025 (rst, clk, r1024_out, r1025_out);
	reg32 r1026 (rst, clk, r1025_out, r1026_out);
	reg32 r1027 (rst, clk, r1026_out, r1027_out);
	reg32 r1028 (rst, clk, r1027_out, r1028_out);
	reg32 r1029 (rst, clk, r1028_out, r1029_out);
	reg32 r1030 (rst, clk, r1029_out, r1030_out);
	reg32 r1031 (rst, clk, r1030_out, r1031_out);
	reg32 r1032 (rst, clk, r1031_out, r1032_out);
	reg32 r1033 (rst, clk, r1032_out, r1033_out);
	reg32 r1034 (rst, clk, r1033_out, r1034_out);
	reg32 r1035 (rst, clk, r1034_out, r1035_out);
	reg32 r1036 (rst, clk, r1035_out, r1036_out);
	reg32 r1037 (rst, clk, r1036_out, r1037_out);
	reg32 r1038 (rst, clk, r1037_out, r1038_out);
	reg32 r1039 (rst, clk, r1038_out, r1039_out);
	reg32 r1040 (rst, clk, r1039_out, r1040_out);
	reg32 r1041 (rst, clk, r1040_out, r1041_out);
	reg32 r1042 (rst, clk, r1041_out, r1042_out);
	reg32 r1043 (rst, clk, r1042_out, r1043_out);
	reg32 r1044 (rst, clk, r1043_out, r1044_out);
	reg32 r1045 (rst, clk, r1044_out, r1045_out);
	reg32 r1046 (rst, clk, r1045_out, r1046_out);
	reg32 r1047 (rst, clk, r1046_out, r1047_out);
	reg32 r1048 (rst, clk, r1047_out, r1048_out);
	reg32 r1049 (rst, clk, r1048_out, r1049_out);
	reg32 r1050 (rst, clk, r1049_out, r1050_out);
	reg32 r1051 (rst, clk, r1050_out, r1051_out);
	reg32 r1052 (rst, clk, r1051_out, r1052_out);
	reg32 r1053 (rst, clk, r1052_out, r1053_out);
	reg32 r1054 (rst, clk, r1053_out, r1054_out);
	reg32 r1055 (rst, clk, r1054_out, r1055_out);
	reg32 r1056 (rst, clk, r1055_out, r1056_out);
	reg32 r1057 (rst, clk, r1056_out, r1057_out);
	reg32 r1058 (rst, clk, r1057_out, r1058_out);
	reg32 r1059 (rst, clk, r1058_out, r1059_out);
	reg32 r1060 (rst, clk, r1059_out, r1060_out);
	reg32 r1061 (rst, clk, r1060_out, r1061_out);
	reg32 r1062 (rst, clk, r1061_out, r1062_out);
	reg32 r1063 (rst, clk, r1062_out, r1063_out);
	reg32 r1064 (rst, clk, r1063_out, r1064_out);
	reg32 r1065 (rst, clk, r1064_out, r1065_out);
	reg32 r1066 (rst, clk, r1065_out, r1066_out);
	reg32 r1067 (rst, clk, r1066_out, r1067_out);
	reg32 r1068 (rst, clk, r1067_out, r1068_out);
	reg32 r1069 (rst, clk, r1068_out, r1069_out);
	reg32 r1070 (rst, clk, r1069_out, r1070_out);
	reg32 r1071 (rst, clk, r1070_out, r1071_out);
	reg32 r1072 (rst, clk, r1071_out, r1072_out);
	reg32 r1073 (rst, clk, r1072_out, r1073_out);
	reg32 r1074 (rst, clk, r1073_out, r1074_out);
	reg32 r1075 (rst, clk, r1074_out, r1075_out);
	reg32 r1076 (rst, clk, r1075_out, r1076_out);
	reg32 r1077 (rst, clk, r1076_out, r1077_out);
	reg32 r1078 (rst, clk, r1077_out, r1078_out);
	reg32 r1079 (rst, clk, r1078_out, r1079_out);
	reg32 r1080 (rst, clk, r1079_out, r1080_out);
	reg32 r1081 (rst, clk, r1080_out, r1081_out);
	reg32 r1082 (rst, clk, r1081_out, r1082_out);
	reg32 r1083 (rst, clk, r1082_out, r1083_out);
	reg32 r1084 (rst, clk, r1083_out, r1084_out);
	reg32 r1085 (rst, clk, r1084_out, r1085_out);
	reg32 r1086 (rst, clk, r1085_out, r1086_out);
	reg32 r1087 (rst, clk, r1086_out, r1087_out);
	reg32 r1088 (rst, clk, r1087_out, r1088_out);
	reg32 r1089 (rst, clk, r1088_out, r1089_out);
	reg32 r1090 (rst, clk, r1089_out, r1090_out);
	reg32 r1091 (rst, clk, r1090_out, r1091_out);
	reg32 r1092 (rst, clk, r1091_out, r1092_out);
	reg32 r1093 (rst, clk, r1092_out, r1093_out);
	reg32 r1094 (rst, clk, r1093_out, r1094_out);
	reg32 r1095 (rst, clk, r1094_out, r1095_out);
	reg32 r1096 (rst, clk, r1095_out, r1096_out);
	reg32 r1097 (rst, clk, r1096_out, r1097_out);
	reg32 r1098 (rst, clk, r1097_out, r1098_out);
	reg32 r1099 (rst, clk, r1098_out, r1099_out);
	reg32 r1100 (rst, clk, r1099_out, r1100_out);
	reg32 r1101 (rst, clk, r1100_out, r1101_out);
	reg32 r1102 (rst, clk, r1101_out, r1102_out);
	reg32 r1103 (rst, clk, r1102_out, r1103_out);
	reg32 r1104 (rst, clk, r1103_out, r1104_out);
	reg32 r1105 (rst, clk, r1104_out, r1105_out);
	reg32 r1106 (rst, clk, r1105_out, r1106_out);
	reg32 r1107 (rst, clk, r1106_out, r1107_out);
	reg32 r1108 (rst, clk, r1107_out, r1108_out);
	reg32 r1109 (rst, clk, r1108_out, r1109_out);
	reg32 r1110 (rst, clk, r1109_out, r1110_out);
	reg32 r1111 (rst, clk, r1110_out, r1111_out);
	reg32 r1112 (rst, clk, r1111_out, r1112_out);
	reg32 r1113 (rst, clk, r1112_out, r1113_out);
	reg32 r1114 (rst, clk, r1113_out, r1114_out);
	reg32 r1115 (rst, clk, r1114_out, r1115_out);
	reg32 r1116 (rst, clk, r1115_out, r1116_out);
	reg32 r1117 (rst, clk, r1116_out, r1117_out);
	reg32 r1118 (rst, clk, r1117_out, r1118_out);
	reg32 r1119 (rst, clk, r1118_out, r1119_out);
	reg32 r1120 (rst, clk, r1119_out, r1120_out);
	reg32 r1121 (rst, clk, r1120_out, r1121_out);
	reg32 r1122 (rst, clk, r1121_out, r1122_out);
	reg32 r1123 (rst, clk, r1122_out, r1123_out);
	reg32 r1124 (rst, clk, r1123_out, r1124_out);
	reg32 r1125 (rst, clk, r1124_out, r1125_out);
	reg32 r1126 (rst, clk, r1125_out, r1126_out);
	reg32 r1127 (rst, clk, r1126_out, r1127_out);
	reg32 r1128 (rst, clk, r1127_out, r1128_out);
	reg32 r1129 (rst, clk, r1128_out, r1129_out);
	reg32 r1130 (rst, clk, r1129_out, r1130_out);
	reg32 r1131 (rst, clk, r1130_out, r1131_out);
	reg32 r1132 (rst, clk, r1131_out, r1132_out);
	reg32 r1133 (rst, clk, r1132_out, r1133_out);
	reg32 r1134 (rst, clk, r1133_out, r1134_out);
	reg32 r1135 (rst, clk, r1134_out, r1135_out);
	reg32 r1136 (rst, clk, r1135_out, r1136_out);
	reg32 r1137 (rst, clk, r1136_out, r1137_out);
	reg32 r1138 (rst, clk, r1137_out, r1138_out);
	reg32 r1139 (rst, clk, r1138_out, r1139_out);
	reg32 r1140 (rst, clk, r1139_out, r1140_out);
	reg32 r1141 (rst, clk, r1140_out, r1141_out);
	reg32 r1142 (rst, clk, r1141_out, r1142_out);
	reg32 r1143 (rst, clk, r1142_out, r1143_out);
	reg32 r1144 (rst, clk, r1143_out, r1144_out);
	reg32 r1145 (rst, clk, r1144_out, r1145_out);
	reg32 r1146 (rst, clk, r1145_out, r1146_out);
	reg32 r1147 (rst, clk, r1146_out, r1147_out);
	reg32 r1148 (rst, clk, r1147_out, r1148_out);
	reg32 r1149 (rst, clk, r1148_out, r1149_out);
	reg32 r1150 (rst, clk, r1149_out, r1150_out);
	reg32 r1151 (rst, clk, r1150_out, r1151_out);
	reg32 r1152 (rst, clk, r1151_out, r1152_out);
	reg32 r1153 (rst, clk, r1152_out, r1153_out);
	reg32 r1154 (rst, clk, r1153_out, r1154_out);
	reg32 r1155 (rst, clk, r1154_out, r1155_out);
	reg32 r1156 (rst, clk, r1155_out, r1156_out);
	reg32 r1157 (rst, clk, r1156_out, r1157_out);
	reg32 r1158 (rst, clk, r1157_out, r1158_out);
	reg32 r1159 (rst, clk, r1158_out, r1159_out);
	reg32 r1160 (rst, clk, r1159_out, r1160_out);
	reg32 r1161 (rst, clk, r1160_out, r1161_out);
	reg32 r1162 (rst, clk, r1161_out, r1162_out);
	reg32 r1163 (rst, clk, r1162_out, r1163_out);
	reg32 r1164 (rst, clk, r1163_out, r1164_out);
	reg32 r1165 (rst, clk, r1164_out, r1165_out);
	reg32 r1166 (rst, clk, r1165_out, r1166_out);
	reg32 r1167 (rst, clk, r1166_out, r1167_out);
	reg32 r1168 (rst, clk, r1167_out, r1168_out);
	reg32 r1169 (rst, clk, r1168_out, r1169_out);
	reg32 r1170 (rst, clk, r1169_out, r1170_out);
	reg32 r1171 (rst, clk, r1170_out, r1171_out);
	reg32 r1172 (rst, clk, r1171_out, r1172_out);
	reg32 r1173 (rst, clk, r1172_out, r1173_out);
	reg32 r1174 (rst, clk, r1173_out, r1174_out);
	reg32 r1175 (rst, clk, r1174_out, r1175_out);
	reg32 r1176 (rst, clk, r1175_out, r1176_out);
	reg32 r1177 (rst, clk, r1176_out, r1177_out);
	reg32 r1178 (rst, clk, r1177_out, r1178_out);
	reg32 r1179 (rst, clk, r1178_out, r1179_out);
	reg32 r1180 (rst, clk, r1179_out, r1180_out);
	reg32 r1181 (rst, clk, r1180_out, r1181_out);
	reg32 r1182 (rst, clk, r1181_out, r1182_out);
	reg32 r1183 (rst, clk, r1182_out, r1183_out);
	reg32 r1184 (rst, clk, r1183_out, r1184_out);
	reg32 r1185 (rst, clk, r1184_out, r1185_out);
	reg32 r1186 (rst, clk, r1185_out, r1186_out);
	reg32 r1187 (rst, clk, r1186_out, r1187_out);
	reg32 r1188 (rst, clk, r1187_out, r1188_out);
	reg32 r1189 (rst, clk, r1188_out, r1189_out);
	reg32 r1190 (rst, clk, r1189_out, r1190_out);
	reg32 r1191 (rst, clk, r1190_out, r1191_out);
	reg32 r1192 (rst, clk, r1191_out, r1192_out);
	reg32 r1193 (rst, clk, r1192_out, r1193_out);
	reg32 r1194 (rst, clk, r1193_out, r1194_out);
	reg32 r1195 (rst, clk, r1194_out, r1195_out);
	reg32 r1196 (rst, clk, r1195_out, r1196_out);
	reg32 r1197 (rst, clk, r1196_out, r1197_out);
	reg32 r1198 (rst, clk, r1197_out, r1198_out);
	reg32 r1199 (rst, clk, r1198_out, r1199_out);
	reg32 r1200 (rst, clk, r1199_out, r1200_out);
	reg32 r1201 (rst, clk, r1200_out, r1201_out);
	reg32 r1202 (rst, clk, r1201_out, r1202_out);
	reg32 r1203 (rst, clk, r1202_out, r1203_out);
	reg32 r1204 (rst, clk, r1203_out, r1204_out);
	reg32 r1205 (rst, clk, r1204_out, r1205_out);
	reg32 r1206 (rst, clk, r1205_out, r1206_out);
	reg32 r1207 (rst, clk, r1206_out, r1207_out);
	reg32 r1208 (rst, clk, r1207_out, r1208_out);
	reg32 r1209 (rst, clk, r1208_out, r1209_out);
	reg32 r1210 (rst, clk, r1209_out, r1210_out);
	reg32 r1211 (rst, clk, r1210_out, r1211_out);
	reg32 r1212 (rst, clk, r1211_out, r1212_out);
	reg32 r1213 (rst, clk, r1212_out, r1213_out);
	reg32 r1214 (rst, clk, r1213_out, r1214_out);
	reg32 r1215 (rst, clk, r1214_out, r1215_out);
	reg32 r1216 (rst, clk, r1215_out, r1216_out);
	reg32 r1217 (rst, clk, r1216_out, r1217_out);
	reg32 r1218 (rst, clk, r1217_out, r1218_out);
	reg32 r1219 (rst, clk, r1218_out, r1219_out);
	reg32 r1220 (rst, clk, r1219_out, r1220_out);
	reg32 r1221 (rst, clk, r1220_out, r1221_out);
	reg32 r1222 (rst, clk, r1221_out, r1222_out);
	reg32 r1223 (rst, clk, r1222_out, r1223_out);
	reg32 r1224 (rst, clk, r1223_out, r1224_out);
	reg32 r1225 (rst, clk, r1224_out, r1225_out);
	reg32 r1226 (rst, clk, r1225_out, r1226_out);
	reg32 r1227 (rst, clk, r1226_out, r1227_out);
	reg32 r1228 (rst, clk, r1227_out, r1228_out);
	reg32 r1229 (rst, clk, r1228_out, r1229_out);
	reg32 r1230 (rst, clk, r1229_out, r1230_out);
	reg32 r1231 (rst, clk, r1230_out, r1231_out);
	reg32 r1232 (rst, clk, r1231_out, r1232_out);
	reg32 r1233 (rst, clk, r1232_out, r1233_out);
	reg32 r1234 (rst, clk, r1233_out, r1234_out);
	reg32 r1235 (rst, clk, r1234_out, r1235_out);
	reg32 r1236 (rst, clk, r1235_out, r1236_out);
	reg32 r1237 (rst, clk, r1236_out, r1237_out);
	reg32 r1238 (rst, clk, r1237_out, r1238_out);
	reg32 r1239 (rst, clk, r1238_out, r1239_out);
	reg32 r1240 (rst, clk, r1239_out, r1240_out);
	reg32 r1241 (rst, clk, r1240_out, r1241_out);
	reg32 r1242 (rst, clk, r1241_out, r1242_out);
	reg32 r1243 (rst, clk, r1242_out, r1243_out);
	reg32 r1244 (rst, clk, r1243_out, r1244_out);
	reg32 r1245 (rst, clk, r1244_out, r1245_out);
	reg32 r1246 (rst, clk, r1245_out, r1246_out);
	reg32 r1247 (rst, clk, r1246_out, r1247_out);
	reg32 r1248 (rst, clk, r1247_out, r1248_out);
	reg32 r1249 (rst, clk, r1248_out, r1249_out);
	reg32 r1250 (rst, clk, r1249_out, r1250_out);
	reg32 r1251 (rst, clk, r1250_out, r1251_out);
	reg32 r1252 (rst, clk, r1251_out, r1252_out);
	reg32 r1253 (rst, clk, r1252_out, r1253_out);
	reg32 r1254 (rst, clk, r1253_out, r1254_out);
	reg32 r1255 (rst, clk, r1254_out, r1255_out);
	reg32 r1256 (rst, clk, r1255_out, r1256_out);
	reg32 r1257 (rst, clk, r1256_out, r1257_out);
	reg32 r1258 (rst, clk, r1257_out, r1258_out);
	reg32 r1259 (rst, clk, r1258_out, r1259_out);
	reg32 r1260 (rst, clk, r1259_out, r1260_out);
	reg32 r1261 (rst, clk, r1260_out, r1261_out);
	reg32 r1262 (rst, clk, r1261_out, r1262_out);
	reg32 r1263 (rst, clk, r1262_out, r1263_out);
	reg32 r1264 (rst, clk, r1263_out, r1264_out);
	reg32 r1265 (rst, clk, r1264_out, r1265_out);
	reg32 r1266 (rst, clk, r1265_out, r1266_out);
	reg32 r1267 (rst, clk, r1266_out, r1267_out);
	reg32 r1268 (rst, clk, r1267_out, r1268_out);
	reg32 r1269 (rst, clk, r1268_out, r1269_out);
	reg32 r1270 (rst, clk, r1269_out, r1270_out);
	reg32 r1271 (rst, clk, r1270_out, r1271_out);
	reg32 r1272 (rst, clk, r1271_out, r1272_out);
	reg32 r1273 (rst, clk, r1272_out, r1273_out);
	reg32 r1274 (rst, clk, r1273_out, r1274_out);
	reg32 r1275 (rst, clk, r1274_out, r1275_out);
	reg32 r1276 (rst, clk, r1275_out, r1276_out);
	reg32 r1277 (rst, clk, r1276_out, r1277_out);
	reg32 r1278 (rst, clk, r1277_out, r1278_out);
	reg32 r1279 (rst, clk, r1278_out, r1279_out);
	reg32 r1280 (rst, clk, r1279_out, r1280_out);
	reg32 r1281 (rst, clk, r1280_out, r1281_out);
	reg32 r1282 (rst, clk, r1281_out, r1282_out);
	reg32 r1283 (rst, clk, r1282_out, r1283_out);
	reg32 r1284 (rst, clk, r1283_out, r1284_out);
	reg32 r1285 (rst, clk, r1284_out, r1285_out);
	reg32 r1286 (rst, clk, r1285_out, r1286_out);
	reg32 r1287 (rst, clk, r1286_out, r1287_out);
	reg32 r1288 (rst, clk, r1287_out, r1288_out);
	reg32 r1289 (rst, clk, r1288_out, r1289_out);
	reg32 r1290 (rst, clk, r1289_out, r1290_out);
	reg32 r1291 (rst, clk, r1290_out, r1291_out);
	reg32 r1292 (rst, clk, r1291_out, r1292_out);
	reg32 r1293 (rst, clk, r1292_out, r1293_out);
	reg32 r1294 (rst, clk, r1293_out, r1294_out);
	reg32 r1295 (rst, clk, r1294_out, r1295_out);
	reg32 r1296 (rst, clk, r1295_out, r1296_out);
	reg32 r1297 (rst, clk, r1296_out, r1297_out);
	reg32 r1298 (rst, clk, r1297_out, r1298_out);
	reg32 r1299 (rst, clk, r1298_out, r1299_out);
	reg32 r1300 (rst, clk, r1299_out, r1300_out);
	reg32 r1301 (rst, clk, r1300_out, r1301_out);
	reg32 r1302 (rst, clk, r1301_out, r1302_out);
	reg32 r1303 (rst, clk, r1302_out, r1303_out);
	reg32 r1304 (rst, clk, r1303_out, r1304_out);
	reg32 r1305 (rst, clk, r1304_out, r1305_out);
	reg32 r1306 (rst, clk, r1305_out, r1306_out);
	reg32 r1307 (rst, clk, r1306_out, r1307_out);
	reg32 r1308 (rst, clk, r1307_out, r1308_out);
	reg32 r1309 (rst, clk, r1308_out, r1309_out);
	reg32 r1310 (rst, clk, r1309_out, r1310_out);
	reg32 r1311 (rst, clk, r1310_out, r1311_out);
	reg32 r1312 (rst, clk, r1311_out, r1312_out);
	reg32 r1313 (rst, clk, r1312_out, r1313_out);
	reg32 r1314 (rst, clk, r1313_out, r1314_out);
	reg32 r1315 (rst, clk, r1314_out, r1315_out);
	reg32 r1316 (rst, clk, r1315_out, r1316_out);
	reg32 r1317 (rst, clk, r1316_out, r1317_out);
	reg32 r1318 (rst, clk, r1317_out, r1318_out);
	reg32 r1319 (rst, clk, r1318_out, r1319_out);
	reg32 r1320 (rst, clk, r1319_out, r1320_out);
	reg32 r1321 (rst, clk, r1320_out, r1321_out);
	reg32 r1322 (rst, clk, r1321_out, r1322_out);
	reg32 r1323 (rst, clk, r1322_out, r1323_out);
	reg32 r1324 (rst, clk, r1323_out, r1324_out);
	reg32 r1325 (rst, clk, r1324_out, r1325_out);
	reg32 r1326 (rst, clk, r1325_out, r1326_out);
	reg32 r1327 (rst, clk, r1326_out, r1327_out);
	reg32 r1328 (rst, clk, r1327_out, r1328_out);
	reg32 r1329 (rst, clk, r1328_out, r1329_out);
	reg32 r1330 (rst, clk, r1329_out, r1330_out);
	reg32 r1331 (rst, clk, r1330_out, r1331_out);
	reg32 r1332 (rst, clk, r1331_out, r1332_out);
	reg32 r1333 (rst, clk, r1332_out, r1333_out);
	reg32 r1334 (rst, clk, r1333_out, r1334_out);
	reg32 r1335 (rst, clk, r1334_out, r1335_out);
	reg32 r1336 (rst, clk, r1335_out, r1336_out);
	reg32 r1337 (rst, clk, r1336_out, r1337_out);
	reg32 r1338 (rst, clk, r1337_out, r1338_out);
	reg32 r1339 (rst, clk, r1338_out, r1339_out);
	reg32 r1340 (rst, clk, r1339_out, r1340_out);
	reg32 r1341 (rst, clk, r1340_out, r1341_out);
	reg32 r1342 (rst, clk, r1341_out, r1342_out);
	reg32 r1343 (rst, clk, r1342_out, r1343_out);
	reg32 r1344 (rst, clk, r1343_out, r1344_out);
	reg32 r1345 (rst, clk, r1344_out, r1345_out);
	reg32 r1346 (rst, clk, r1345_out, r1346_out);
	reg32 r1347 (rst, clk, r1346_out, r1347_out);
	reg32 r1348 (rst, clk, r1347_out, r1348_out);
	reg32 r1349 (rst, clk, r1348_out, r1349_out);
	reg32 r1350 (rst, clk, r1349_out, r1350_out);
	reg32 r1351 (rst, clk, r1350_out, r1351_out);
	reg32 r1352 (rst, clk, r1351_out, r1352_out);
	reg32 r1353 (rst, clk, r1352_out, r1353_out);
	reg32 r1354 (rst, clk, r1353_out, r1354_out);
	reg32 r1355 (rst, clk, r1354_out, r1355_out);
	reg32 r1356 (rst, clk, r1355_out, r1356_out);
	reg32 r1357 (rst, clk, r1356_out, r1357_out);
	reg32 r1358 (rst, clk, r1357_out, r1358_out);
	reg32 r1359 (rst, clk, r1358_out, r1359_out);
	reg32 r1360 (rst, clk, r1359_out, r1360_out);
	reg32 r1361 (rst, clk, r1360_out, r1361_out);
	reg32 r1362 (rst, clk, r1361_out, r1362_out);
	reg32 r1363 (rst, clk, r1362_out, r1363_out);
	reg32 r1364 (rst, clk, r1363_out, r1364_out);
	reg32 r1365 (rst, clk, r1364_out, r1365_out);
	reg32 r1366 (rst, clk, r1365_out, r1366_out);
	reg32 r1367 (rst, clk, r1366_out, r1367_out);
	reg32 r1368 (rst, clk, r1367_out, r1368_out);
	reg32 r1369 (rst, clk, r1368_out, r1369_out);
	reg32 r1370 (rst, clk, r1369_out, r1370_out);
	reg32 r1371 (rst, clk, r1370_out, r1371_out);
	reg32 r1372 (rst, clk, r1371_out, r1372_out);
	reg32 r1373 (rst, clk, r1372_out, r1373_out);
	reg32 r1374 (rst, clk, r1373_out, r1374_out);
	reg32 r1375 (rst, clk, r1374_out, r1375_out);
	reg32 r1376 (rst, clk, r1375_out, r1376_out);
	reg32 r1377 (rst, clk, r1376_out, r1377_out);
	reg32 r1378 (rst, clk, r1377_out, r1378_out);
	reg32 r1379 (rst, clk, r1378_out, r1379_out);
	reg32 r1380 (rst, clk, r1379_out, r1380_out);
	reg32 r1381 (rst, clk, r1380_out, r1381_out);
	reg32 r1382 (rst, clk, r1381_out, r1382_out);
	reg32 r1383 (rst, clk, r1382_out, r1383_out);
	reg32 r1384 (rst, clk, r1383_out, r1384_out);
	reg32 r1385 (rst, clk, r1384_out, r1385_out);
	reg32 r1386 (rst, clk, r1385_out, r1386_out);
	reg32 r1387 (rst, clk, r1386_out, r1387_out);
	reg32 r1388 (rst, clk, r1387_out, r1388_out);
	reg32 r1389 (rst, clk, r1388_out, r1389_out);
	reg32 r1390 (rst, clk, r1389_out, r1390_out);
	reg32 r1391 (rst, clk, r1390_out, r1391_out);
	reg32 r1392 (rst, clk, r1391_out, r1392_out);
	reg32 r1393 (rst, clk, r1392_out, r1393_out);
	reg32 r1394 (rst, clk, r1393_out, r1394_out);
	reg32 r1395 (rst, clk, r1394_out, r1395_out);
	reg32 r1396 (rst, clk, r1395_out, r1396_out);
	reg32 r1397 (rst, clk, r1396_out, r1397_out);
	reg32 r1398 (rst, clk, r1397_out, r1398_out);
	reg32 r1399 (rst, clk, r1398_out, r1399_out);
	reg32 r1400 (rst, clk, r1399_out, r1400_out);
	reg32 r1401 (rst, clk, r1400_out, r1401_out);
	reg32 r1402 (rst, clk, r1401_out, r1402_out);
	reg32 r1403 (rst, clk, r1402_out, r1403_out);
	reg32 r1404 (rst, clk, r1403_out, r1404_out);
	reg32 r1405 (rst, clk, r1404_out, r1405_out);
	reg32 r1406 (rst, clk, r1405_out, r1406_out);
	reg32 r1407 (rst, clk, r1406_out, r1407_out);
	reg32 r1408 (rst, clk, r1407_out, r1408_out);
	reg32 r1409 (rst, clk, r1408_out, r1409_out);
	reg32 r1410 (rst, clk, r1409_out, r1410_out);
	reg32 r1411 (rst, clk, r1410_out, r1411_out);
	reg32 r1412 (rst, clk, r1411_out, r1412_out);
	reg32 r1413 (rst, clk, r1412_out, r1413_out);
	reg32 r1414 (rst, clk, r1413_out, r1414_out);
	reg32 r1415 (rst, clk, r1414_out, r1415_out);
	reg32 r1416 (rst, clk, r1415_out, r1416_out);
	reg32 r1417 (rst, clk, r1416_out, r1417_out);
	reg32 r1418 (rst, clk, r1417_out, r1418_out);
	reg32 r1419 (rst, clk, r1418_out, r1419_out);
	reg32 r1420 (rst, clk, r1419_out, r1420_out);
	reg32 r1421 (rst, clk, r1420_out, r1421_out);
	reg32 r1422 (rst, clk, r1421_out, r1422_out);
	reg32 r1423 (rst, clk, r1422_out, r1423_out);
	reg32 r1424 (rst, clk, r1423_out, r1424_out);
	reg32 r1425 (rst, clk, r1424_out, r1425_out);
	reg32 r1426 (rst, clk, r1425_out, r1426_out);
	reg32 r1427 (rst, clk, r1426_out, r1427_out);
	reg32 r1428 (rst, clk, r1427_out, r1428_out);
	reg32 r1429 (rst, clk, r1428_out, r1429_out);
	reg32 r1430 (rst, clk, r1429_out, r1430_out);
	reg32 r1431 (rst, clk, r1430_out, r1431_out);
	reg32 r1432 (rst, clk, r1431_out, r1432_out);
	reg32 r1433 (rst, clk, r1432_out, r1433_out);
	reg32 r1434 (rst, clk, r1433_out, r1434_out);
	reg32 r1435 (rst, clk, r1434_out, r1435_out);
	reg32 r1436 (rst, clk, r1435_out, r1436_out);
	reg32 r1437 (rst, clk, r1436_out, r1437_out);
	reg32 r1438 (rst, clk, r1437_out, r1438_out);
	reg32 r1439 (rst, clk, r1438_out, r1439_out);
	reg32 r1440 (rst, clk, r1439_out, r1440_out);
	reg32 r1441 (rst, clk, r1440_out, r1441_out);
	reg32 r1442 (rst, clk, r1441_out, r1442_out);
	reg32 r1443 (rst, clk, r1442_out, r1443_out);
	reg32 r1444 (rst, clk, r1443_out, r1444_out);
	reg32 r1445 (rst, clk, r1444_out, r1445_out);
	reg32 r1446 (rst, clk, r1445_out, r1446_out);
	reg32 r1447 (rst, clk, r1446_out, r1447_out);
	reg32 r1448 (rst, clk, r1447_out, r1448_out);
	reg32 r1449 (rst, clk, r1448_out, r1449_out);
	reg32 r1450 (rst, clk, r1449_out, r1450_out);
	reg32 r1451 (rst, clk, r1450_out, r1451_out);
	reg32 r1452 (rst, clk, r1451_out, r1452_out);
	reg32 r1453 (rst, clk, r1452_out, r1453_out);
	reg32 r1454 (rst, clk, r1453_out, r1454_out);
	reg32 r1455 (rst, clk, r1454_out, r1455_out);
	reg32 r1456 (rst, clk, r1455_out, r1456_out);
	reg32 r1457 (rst, clk, r1456_out, r1457_out);
	reg32 r1458 (rst, clk, r1457_out, r1458_out);
	reg32 r1459 (rst, clk, r1458_out, r1459_out);
	reg32 r1460 (rst, clk, r1459_out, r1460_out);
	reg32 r1461 (rst, clk, r1460_out, r1461_out);
	reg32 r1462 (rst, clk, r1461_out, r1462_out);
	reg32 r1463 (rst, clk, r1462_out, r1463_out);
	reg32 r1464 (rst, clk, r1463_out, r1464_out);
	reg32 r1465 (rst, clk, r1464_out, r1465_out);
	reg32 r1466 (rst, clk, r1465_out, r1466_out);
	reg32 r1467 (rst, clk, r1466_out, r1467_out);
	reg32 r1468 (rst, clk, r1467_out, r1468_out);
	reg32 r1469 (rst, clk, r1468_out, r1469_out);
	reg32 r1470 (rst, clk, r1469_out, r1470_out);
	reg32 r1471 (rst, clk, r1470_out, r1471_out);
	reg32 r1472 (rst, clk, r1471_out, r1472_out);
	reg32 r1473 (rst, clk, r1472_out, r1473_out);
	reg32 r1474 (rst, clk, r1473_out, r1474_out);
	reg32 r1475 (rst, clk, r1474_out, r1475_out);
	reg32 r1476 (rst, clk, r1475_out, r1476_out);
	reg32 r1477 (rst, clk, r1476_out, r1477_out);
	reg32 r1478 (rst, clk, r1477_out, r1478_out);
	reg32 r1479 (rst, clk, r1478_out, r1479_out);
	reg32 r1480 (rst, clk, r1479_out, r1480_out);
	reg32 r1481 (rst, clk, r1480_out, r1481_out);
	reg32 r1482 (rst, clk, r1481_out, r1482_out);
	reg32 r1483 (rst, clk, r1482_out, r1483_out);
	reg32 r1484 (rst, clk, r1483_out, r1484_out);
	reg32 r1485 (rst, clk, r1484_out, r1485_out);
	reg32 r1486 (rst, clk, r1485_out, r1486_out);
	reg32 r1487 (rst, clk, r1486_out, r1487_out);
	reg32 r1488 (rst, clk, r1487_out, r1488_out);
	reg32 r1489 (rst, clk, r1488_out, r1489_out);
	reg32 r1490 (rst, clk, r1489_out, r1490_out);
	reg32 r1491 (rst, clk, r1490_out, r1491_out);
	reg32 r1492 (rst, clk, r1491_out, r1492_out);
	reg32 r1493 (rst, clk, r1492_out, r1493_out);
	reg32 r1494 (rst, clk, r1493_out, r1494_out);
	reg32 r1495 (rst, clk, r1494_out, r1495_out);
	reg32 r1496 (rst, clk, r1495_out, r1496_out);
	reg32 r1497 (rst, clk, r1496_out, r1497_out);
	reg32 r1498 (rst, clk, r1497_out, r1498_out);
	reg32 r1499 (rst, clk, r1498_out, r1499_out);
	reg32 r1500 (rst, clk, r1499_out, r1500_out);
	reg32 r1501 (rst, clk, r1500_out, r1501_out);
	reg32 r1502 (rst, clk, r1501_out, r1502_out);
	reg32 r1503 (rst, clk, r1502_out, r1503_out);
	reg32 r1504 (rst, clk, r1503_out, r1504_out);
	reg32 r1505 (rst, clk, r1504_out, r1505_out);
	reg32 r1506 (rst, clk, r1505_out, r1506_out);
	reg32 r1507 (rst, clk, r1506_out, r1507_out);
	reg32 r1508 (rst, clk, r1507_out, r1508_out);
	reg32 r1509 (rst, clk, r1508_out, r1509_out);
	reg32 r1510 (rst, clk, r1509_out, r1510_out);
	reg32 r1511 (rst, clk, r1510_out, r1511_out);
	reg32 r1512 (rst, clk, r1511_out, r1512_out);
	reg32 r1513 (rst, clk, r1512_out, r1513_out);
	reg32 r1514 (rst, clk, r1513_out, r1514_out);
	reg32 r1515 (rst, clk, r1514_out, r1515_out);
	reg32 r1516 (rst, clk, r1515_out, r1516_out);
	reg32 r1517 (rst, clk, r1516_out, r1517_out);
	reg32 r1518 (rst, clk, r1517_out, r1518_out);
	reg32 r1519 (rst, clk, r1518_out, r1519_out);
	reg32 r1520 (rst, clk, r1519_out, r1520_out);
	reg32 r1521 (rst, clk, r1520_out, r1521_out);
	reg32 r1522 (rst, clk, r1521_out, r1522_out);
	reg32 r1523 (rst, clk, r1522_out, r1523_out);
	reg32 r1524 (rst, clk, r1523_out, r1524_out);
	reg32 r1525 (rst, clk, r1524_out, r1525_out);
	reg32 r1526 (rst, clk, r1525_out, r1526_out);
	reg32 r1527 (rst, clk, r1526_out, r1527_out);
	reg32 r1528 (rst, clk, r1527_out, r1528_out);
	reg32 r1529 (rst, clk, r1528_out, r1529_out);
	reg32 r1530 (rst, clk, r1529_out, r1530_out);
	reg32 r1531 (rst, clk, r1530_out, r1531_out);
	reg32 r1532 (rst, clk, r1531_out, r1532_out);
	reg32 r1533 (rst, clk, r1532_out, r1533_out);
	reg32 r1534 (rst, clk, r1533_out, r1534_out);
	reg32 r1535 (rst, clk, r1534_out, r1535_out);
	reg32 r1536 (rst, clk, r1535_out, r1536_out);
	reg32 r1537 (rst, clk, r1536_out, r1537_out);
	reg32 r1538 (rst, clk, r1537_out, r1538_out);
	reg32 r1539 (rst, clk, r1538_out, r1539_out);
	reg32 r1540 (rst, clk, r1539_out, r1540_out);
	reg32 r1541 (rst, clk, r1540_out, r1541_out);
	reg32 r1542 (rst, clk, r1541_out, r1542_out);
	reg32 r1543 (rst, clk, r1542_out, r1543_out);
	reg32 r1544 (rst, clk, r1543_out, r1544_out);
	reg32 r1545 (rst, clk, r1544_out, r1545_out);
	reg32 r1546 (rst, clk, r1545_out, r1546_out);
	reg32 r1547 (rst, clk, r1546_out, r1547_out);
	reg32 r1548 (rst, clk, r1547_out, r1548_out);
	reg32 r1549 (rst, clk, r1548_out, r1549_out);
	reg32 r1550 (rst, clk, r1549_out, r1550_out);
	reg32 r1551 (rst, clk, r1550_out, r1551_out);
	reg32 r1552 (rst, clk, r1551_out, r1552_out);
	reg32 r1553 (rst, clk, r1552_out, r1553_out);
	reg32 r1554 (rst, clk, r1553_out, r1554_out);
	reg32 r1555 (rst, clk, r1554_out, r1555_out);
	reg32 r1556 (rst, clk, r1555_out, r1556_out);
	reg32 r1557 (rst, clk, r1556_out, r1557_out);
	reg32 r1558 (rst, clk, r1557_out, r1558_out);
	reg32 r1559 (rst, clk, r1558_out, r1559_out);
	reg32 r1560 (rst, clk, r1559_out, r1560_out);
	reg32 r1561 (rst, clk, r1560_out, r1561_out);
	reg32 r1562 (rst, clk, r1561_out, r1562_out);
	reg32 r1563 (rst, clk, r1562_out, r1563_out);
	reg32 r1564 (rst, clk, r1563_out, r1564_out);
	reg32 r1565 (rst, clk, r1564_out, r1565_out);
	reg32 r1566 (rst, clk, r1565_out, r1566_out);
	reg32 r1567 (rst, clk, r1566_out, r1567_out);
	reg32 r1568 (rst, clk, r1567_out, r1568_out);
	reg32 r1569 (rst, clk, r1568_out, r1569_out);
	reg32 r1570 (rst, clk, r1569_out, r1570_out);
	reg32 r1571 (rst, clk, r1570_out, r1571_out);
	reg32 r1572 (rst, clk, r1571_out, r1572_out);
	reg32 r1573 (rst, clk, r1572_out, r1573_out);
	reg32 r1574 (rst, clk, r1573_out, r1574_out);
	reg32 r1575 (rst, clk, r1574_out, r1575_out);
	reg32 r1576 (rst, clk, r1575_out, r1576_out);
	reg32 r1577 (rst, clk, r1576_out, r1577_out);
	reg32 r1578 (rst, clk, r1577_out, r1578_out);
	reg32 r1579 (rst, clk, r1578_out, r1579_out);
	reg32 r1580 (rst, clk, r1579_out, r1580_out);
	reg32 r1581 (rst, clk, r1580_out, r1581_out);
	reg32 r1582 (rst, clk, r1581_out, r1582_out);
	reg32 r1583 (rst, clk, r1582_out, r1583_out);
	reg32 r1584 (rst, clk, r1583_out, r1584_out);
	reg32 r1585 (rst, clk, r1584_out, r1585_out);
	reg32 r1586 (rst, clk, r1585_out, r1586_out);
	reg32 r1587 (rst, clk, r1586_out, r1587_out);
	reg32 r1588 (rst, clk, r1587_out, r1588_out);
	reg32 r1589 (rst, clk, r1588_out, r1589_out);
	reg32 r1590 (rst, clk, r1589_out, r1590_out);
	reg32 r1591 (rst, clk, r1590_out, r1591_out);
	reg32 r1592 (rst, clk, r1591_out, r1592_out);
	reg32 r1593 (rst, clk, r1592_out, r1593_out);
	reg32 r1594 (rst, clk, r1593_out, r1594_out);
	reg32 r1595 (rst, clk, r1594_out, r1595_out);
	reg32 r1596 (rst, clk, r1595_out, r1596_out);
	reg32 r1597 (rst, clk, r1596_out, r1597_out);
	reg32 r1598 (rst, clk, r1597_out, r1598_out);
	reg32 r1599 (rst, clk, r1598_out, r1599_out);
	reg32 r1600 (rst, clk, r1599_out, r1600_out);
	reg32 r1601 (rst, clk, r1600_out, r1601_out);
	reg32 r1602 (rst, clk, r1601_out, r1602_out);
	reg32 r1603 (rst, clk, r1602_out, r1603_out);
	reg32 r1604 (rst, clk, r1603_out, r1604_out);
	reg32 r1605 (rst, clk, r1604_out, r1605_out);
	reg32 r1606 (rst, clk, r1605_out, r1606_out);
	reg32 r1607 (rst, clk, r1606_out, r1607_out);
	reg32 r1608 (rst, clk, r1607_out, r1608_out);
	reg32 r1609 (rst, clk, r1608_out, r1609_out);
	reg32 r1610 (rst, clk, r1609_out, r1610_out);
	reg32 r1611 (rst, clk, r1610_out, r1611_out);
	reg32 r1612 (rst, clk, r1611_out, r1612_out);
	reg32 r1613 (rst, clk, r1612_out, r1613_out);
	reg32 r1614 (rst, clk, r1613_out, r1614_out);
	reg32 r1615 (rst, clk, r1614_out, r1615_out);
	reg32 r1616 (rst, clk, r1615_out, r1616_out);
	reg32 r1617 (rst, clk, r1616_out, r1617_out);
	reg32 r1618 (rst, clk, r1617_out, r1618_out);
	reg32 r1619 (rst, clk, r1618_out, r1619_out);
	reg32 r1620 (rst, clk, r1619_out, r1620_out);
	reg32 r1621 (rst, clk, r1620_out, r1621_out);
	reg32 r1622 (rst, clk, r1621_out, r1622_out);
	reg32 r1623 (rst, clk, r1622_out, r1623_out);
	reg32 r1624 (rst, clk, r1623_out, r1624_out);
	reg32 r1625 (rst, clk, r1624_out, r1625_out);
	reg32 r1626 (rst, clk, r1625_out, r1626_out);
	reg32 r1627 (rst, clk, r1626_out, r1627_out);
	reg32 r1628 (rst, clk, r1627_out, r1628_out);
	reg32 r1629 (rst, clk, r1628_out, r1629_out);
	reg32 r1630 (rst, clk, r1629_out, r1630_out);
	reg32 r1631 (rst, clk, r1630_out, r1631_out);
	reg32 r1632 (rst, clk, r1631_out, r1632_out);
	reg32 r1633 (rst, clk, r1632_out, r1633_out);
	reg32 r1634 (rst, clk, r1633_out, r1634_out);
	reg32 r1635 (rst, clk, r1634_out, r1635_out);
	reg32 r1636 (rst, clk, r1635_out, r1636_out);
	reg32 r1637 (rst, clk, r1636_out, r1637_out);
	reg32 r1638 (rst, clk, r1637_out, r1638_out);
	reg32 r1639 (rst, clk, r1638_out, r1639_out);
	reg32 r1640 (rst, clk, r1639_out, r1640_out);
	reg32 r1641 (rst, clk, r1640_out, r1641_out);
	reg32 r1642 (rst, clk, r1641_out, r1642_out);
	reg32 r1643 (rst, clk, r1642_out, r1643_out);
	reg32 r1644 (rst, clk, r1643_out, r1644_out);
	reg32 r1645 (rst, clk, r1644_out, r1645_out);
	reg32 r1646 (rst, clk, r1645_out, r1646_out);
	reg32 r1647 (rst, clk, r1646_out, r1647_out);
	reg32 r1648 (rst, clk, r1647_out, r1648_out);
	reg32 r1649 (rst, clk, r1648_out, r1649_out);
	reg32 r1650 (rst, clk, r1649_out, r1650_out);
	reg32 r1651 (rst, clk, r1650_out, r1651_out);
	reg32 r1652 (rst, clk, r1651_out, r1652_out);
	reg32 r1653 (rst, clk, r1652_out, r1653_out);
	reg32 r1654 (rst, clk, r1653_out, r1654_out);
	reg32 r1655 (rst, clk, r1654_out, r1655_out);
	reg32 r1656 (rst, clk, r1655_out, r1656_out);
	reg32 r1657 (rst, clk, r1656_out, r1657_out);
	reg32 r1658 (rst, clk, r1657_out, r1658_out);
	reg32 r1659 (rst, clk, r1658_out, r1659_out);
	reg32 r1660 (rst, clk, r1659_out, r1660_out);
	reg32 r1661 (rst, clk, r1660_out, r1661_out);
	reg32 r1662 (rst, clk, r1661_out, r1662_out);
	reg32 r1663 (rst, clk, r1662_out, r1663_out);
	reg32 r1664 (rst, clk, r1663_out, r1664_out);
	reg32 r1665 (rst, clk, r1664_out, r1665_out);
	reg32 r1666 (rst, clk, r1665_out, r1666_out);
	reg32 r1667 (rst, clk, r1666_out, r1667_out);
	reg32 r1668 (rst, clk, r1667_out, r1668_out);
	reg32 r1669 (rst, clk, r1668_out, r1669_out);
	reg32 r1670 (rst, clk, r1669_out, r1670_out);
	reg32 r1671 (rst, clk, r1670_out, r1671_out);
	reg32 r1672 (rst, clk, r1671_out, r1672_out);
	reg32 r1673 (rst, clk, r1672_out, r1673_out);
	reg32 r1674 (rst, clk, r1673_out, r1674_out);
	reg32 r1675 (rst, clk, r1674_out, r1675_out);
	reg32 r1676 (rst, clk, r1675_out, r1676_out);
	reg32 r1677 (rst, clk, r1676_out, r1677_out);
	reg32 r1678 (rst, clk, r1677_out, r1678_out);
	reg32 r1679 (rst, clk, r1678_out, r1679_out);
	reg32 r1680 (rst, clk, r1679_out, r1680_out);
	reg32 r1681 (rst, clk, r1680_out, r1681_out);
	reg32 r1682 (rst, clk, r1681_out, r1682_out);
	reg32 r1683 (rst, clk, r1682_out, r1683_out);
	reg32 r1684 (rst, clk, r1683_out, r1684_out);
	reg32 r1685 (rst, clk, r1684_out, r1685_out);
	reg32 r1686 (rst, clk, r1685_out, r1686_out);
	reg32 r1687 (rst, clk, r1686_out, r1687_out);
	reg32 r1688 (rst, clk, r1687_out, r1688_out);
	reg32 r1689 (rst, clk, r1688_out, r1689_out);
	reg32 r1690 (rst, clk, r1689_out, r1690_out);
	reg32 r1691 (rst, clk, r1690_out, r1691_out);
	reg32 r1692 (rst, clk, r1691_out, r1692_out);
	reg32 r1693 (rst, clk, r1692_out, r1693_out);
	reg32 r1694 (rst, clk, r1693_out, r1694_out);
	reg32 r1695 (rst, clk, r1694_out, r1695_out);
	reg32 r1696 (rst, clk, r1695_out, r1696_out);
	reg32 r1697 (rst, clk, r1696_out, r1697_out);
	reg32 r1698 (rst, clk, r1697_out, r1698_out);
	reg32 r1699 (rst, clk, r1698_out, r1699_out);
	reg32 r1700 (rst, clk, r1699_out, r1700_out);
	reg32 r1701 (rst, clk, r1700_out, r1701_out);
	reg32 r1702 (rst, clk, r1701_out, r1702_out);
	reg32 r1703 (rst, clk, r1702_out, r1703_out);
	reg32 r1704 (rst, clk, r1703_out, r1704_out);
	reg32 r1705 (rst, clk, r1704_out, r1705_out);
	reg32 r1706 (rst, clk, r1705_out, r1706_out);
	reg32 r1707 (rst, clk, r1706_out, r1707_out);
	reg32 r1708 (rst, clk, r1707_out, r1708_out);
	reg32 r1709 (rst, clk, r1708_out, r1709_out);
	reg32 r1710 (rst, clk, r1709_out, r1710_out);
	reg32 r1711 (rst, clk, r1710_out, r1711_out);
	reg32 r1712 (rst, clk, r1711_out, r1712_out);
	reg32 r1713 (rst, clk, r1712_out, r1713_out);
	reg32 r1714 (rst, clk, r1713_out, r1714_out);
	reg32 r1715 (rst, clk, r1714_out, r1715_out);
	reg32 r1716 (rst, clk, r1715_out, r1716_out);
	reg32 r1717 (rst, clk, r1716_out, r1717_out);
	reg32 r1718 (rst, clk, r1717_out, r1718_out);
	reg32 r1719 (rst, clk, r1718_out, r1719_out);
	reg32 r1720 (rst, clk, r1719_out, r1720_out);
	reg32 r1721 (rst, clk, r1720_out, r1721_out);
	reg32 r1722 (rst, clk, r1721_out, r1722_out);
	reg32 r1723 (rst, clk, r1722_out, r1723_out);
	reg32 r1724 (rst, clk, r1723_out, r1724_out);
	reg32 r1725 (rst, clk, r1724_out, r1725_out);
	reg32 r1726 (rst, clk, r1725_out, r1726_out);
	reg32 r1727 (rst, clk, r1726_out, r1727_out);
	reg32 r1728 (rst, clk, r1727_out, r1728_out);
	reg32 r1729 (rst, clk, r1728_out, r1729_out);
	reg32 r1730 (rst, clk, r1729_out, r1730_out);
	reg32 r1731 (rst, clk, r1730_out, r1731_out);
	reg32 r1732 (rst, clk, r1731_out, r1732_out);
	reg32 r1733 (rst, clk, r1732_out, r1733_out);
	reg32 r1734 (rst, clk, r1733_out, r1734_out);
	reg32 r1735 (rst, clk, r1734_out, r1735_out);
	reg32 r1736 (rst, clk, r1735_out, r1736_out);
	reg32 r1737 (rst, clk, r1736_out, r1737_out);
	reg32 r1738 (rst, clk, r1737_out, r1738_out);
	reg32 r1739 (rst, clk, r1738_out, r1739_out);
	reg32 r1740 (rst, clk, r1739_out, r1740_out);
	reg32 r1741 (rst, clk, r1740_out, r1741_out);
	reg32 r1742 (rst, clk, r1741_out, r1742_out);
	reg32 r1743 (rst, clk, r1742_out, r1743_out);
	reg32 r1744 (rst, clk, r1743_out, r1744_out);
	reg32 r1745 (rst, clk, r1744_out, r1745_out);
	reg32 r1746 (rst, clk, r1745_out, r1746_out);
	reg32 r1747 (rst, clk, r1746_out, r1747_out);
	reg32 r1748 (rst, clk, r1747_out, r1748_out);
	reg32 r1749 (rst, clk, r1748_out, r1749_out);
	reg32 r1750 (rst, clk, r1749_out, r1750_out);
	reg32 r1751 (rst, clk, r1750_out, r1751_out);
	reg32 r1752 (rst, clk, r1751_out, r1752_out);
	reg32 r1753 (rst, clk, r1752_out, r1753_out);
	reg32 r1754 (rst, clk, r1753_out, r1754_out);
	reg32 r1755 (rst, clk, r1754_out, r1755_out);
	reg32 r1756 (rst, clk, r1755_out, r1756_out);
	reg32 r1757 (rst, clk, r1756_out, r1757_out);
	reg32 r1758 (rst, clk, r1757_out, r1758_out);
	reg32 r1759 (rst, clk, r1758_out, r1759_out);
	reg32 r1760 (rst, clk, r1759_out, r1760_out);
	reg32 r1761 (rst, clk, r1760_out, r1761_out);
	reg32 r1762 (rst, clk, r1761_out, r1762_out);
	reg32 r1763 (rst, clk, r1762_out, r1763_out);
	reg32 r1764 (rst, clk, r1763_out, r1764_out);
	reg32 r1765 (rst, clk, r1764_out, r1765_out);
	reg32 r1766 (rst, clk, r1765_out, r1766_out);
	reg32 r1767 (rst, clk, r1766_out, r1767_out);
	reg32 r1768 (rst, clk, r1767_out, r1768_out);
	reg32 r1769 (rst, clk, r1768_out, r1769_out);
	reg32 r1770 (rst, clk, r1769_out, r1770_out);
	reg32 r1771 (rst, clk, r1770_out, r1771_out);
	reg32 r1772 (rst, clk, r1771_out, r1772_out);
	reg32 r1773 (rst, clk, r1772_out, r1773_out);
	reg32 r1774 (rst, clk, r1773_out, r1774_out);
	reg32 r1775 (rst, clk, r1774_out, r1775_out);
	reg32 r1776 (rst, clk, r1775_out, r1776_out);
	reg32 r1777 (rst, clk, r1776_out, r1777_out);
	reg32 r1778 (rst, clk, r1777_out, r1778_out);
	reg32 r1779 (rst, clk, r1778_out, r1779_out);
	reg32 r1780 (rst, clk, r1779_out, r1780_out);
	reg32 r1781 (rst, clk, r1780_out, r1781_out);
	reg32 r1782 (rst, clk, r1781_out, r1782_out);
	reg32 r1783 (rst, clk, r1782_out, r1783_out);
	reg32 r1784 (rst, clk, r1783_out, r1784_out);
	reg32 r1785 (rst, clk, r1784_out, r1785_out);
	reg32 r1786 (rst, clk, r1785_out, r1786_out);
	reg32 r1787 (rst, clk, r1786_out, r1787_out);
	reg32 r1788 (rst, clk, r1787_out, r1788_out);
	reg32 r1789 (rst, clk, r1788_out, r1789_out);
	reg32 r1790 (rst, clk, r1789_out, r1790_out);
	reg32 r1791 (rst, clk, r1790_out, r1791_out);
	reg32 r1792 (rst, clk, r1791_out, r1792_out);
	reg32 r1793 (rst, clk, r1792_out, r1793_out);
	reg32 r1794 (rst, clk, r1793_out, r1794_out);
	reg32 r1795 (rst, clk, r1794_out, r1795_out);
	reg32 r1796 (rst, clk, r1795_out, r1796_out);
	reg32 r1797 (rst, clk, r1796_out, r1797_out);
	reg32 r1798 (rst, clk, r1797_out, r1798_out);
	reg32 r1799 (rst, clk, r1798_out, r1799_out);
	reg32 r1800 (rst, clk, r1799_out, r1800_out);
	reg32 r1801 (rst, clk, r1800_out, r1801_out);
	reg32 r1802 (rst, clk, r1801_out, r1802_out);
	reg32 r1803 (rst, clk, r1802_out, r1803_out);
	reg32 r1804 (rst, clk, r1803_out, r1804_out);
	reg32 r1805 (rst, clk, r1804_out, r1805_out);
	reg32 r1806 (rst, clk, r1805_out, r1806_out);
	reg32 r1807 (rst, clk, r1806_out, r1807_out);
	reg32 r1808 (rst, clk, r1807_out, r1808_out);
	reg32 r1809 (rst, clk, r1808_out, r1809_out);
	reg32 r1810 (rst, clk, r1809_out, r1810_out);
	reg32 r1811 (rst, clk, r1810_out, r1811_out);
	reg32 r1812 (rst, clk, r1811_out, r1812_out);
	reg32 r1813 (rst, clk, r1812_out, r1813_out);
	reg32 r1814 (rst, clk, r1813_out, r1814_out);
	reg32 r1815 (rst, clk, r1814_out, r1815_out);
	reg32 r1816 (rst, clk, r1815_out, r1816_out);
	reg32 r1817 (rst, clk, r1816_out, r1817_out);
	reg32 r1818 (rst, clk, r1817_out, r1818_out);
	reg32 r1819 (rst, clk, r1818_out, r1819_out);
	reg32 r1820 (rst, clk, r1819_out, r1820_out);
	reg32 r1821 (rst, clk, r1820_out, r1821_out);
	reg32 r1822 (rst, clk, r1821_out, r1822_out);
	reg32 r1823 (rst, clk, r1822_out, r1823_out);
	reg32 r1824 (rst, clk, r1823_out, r1824_out);
	reg32 r1825 (rst, clk, r1824_out, r1825_out);
	reg32 r1826 (rst, clk, r1825_out, r1826_out);
	reg32 r1827 (rst, clk, r1826_out, r1827_out);
	reg32 r1828 (rst, clk, r1827_out, r1828_out);
	reg32 r1829 (rst, clk, r1828_out, r1829_out);
	reg32 r1830 (rst, clk, r1829_out, r1830_out);
	reg32 r1831 (rst, clk, r1830_out, r1831_out);
	reg32 r1832 (rst, clk, r1831_out, r1832_out);
	reg32 r1833 (rst, clk, r1832_out, r1833_out);
	reg32 r1834 (rst, clk, r1833_out, r1834_out);
	reg32 r1835 (rst, clk, r1834_out, r1835_out);
	reg32 r1836 (rst, clk, r1835_out, r1836_out);
	reg32 r1837 (rst, clk, r1836_out, r1837_out);
	reg32 r1838 (rst, clk, r1837_out, r1838_out);
	reg32 r1839 (rst, clk, r1838_out, r1839_out);
	reg32 r1840 (rst, clk, r1839_out, r1840_out);
	reg32 r1841 (rst, clk, r1840_out, r1841_out);
	reg32 r1842 (rst, clk, r1841_out, r1842_out);
	reg32 r1843 (rst, clk, r1842_out, r1843_out);
	reg32 r1844 (rst, clk, r1843_out, r1844_out);
	reg32 r1845 (rst, clk, r1844_out, r1845_out);
	reg32 r1846 (rst, clk, r1845_out, r1846_out);
	reg32 r1847 (rst, clk, r1846_out, r1847_out);
	reg32 r1848 (rst, clk, r1847_out, r1848_out);
	reg32 r1849 (rst, clk, r1848_out, r1849_out);
	reg32 r1850 (rst, clk, r1849_out, r1850_out);
	reg32 r1851 (rst, clk, r1850_out, r1851_out);
	reg32 r1852 (rst, clk, r1851_out, r1852_out);
	reg32 r1853 (rst, clk, r1852_out, r1853_out);
	reg32 r1854 (rst, clk, r1853_out, r1854_out);
	reg32 r1855 (rst, clk, r1854_out, r1855_out);
	reg32 r1856 (rst, clk, r1855_out, r1856_out);
	reg32 r1857 (rst, clk, r1856_out, r1857_out);
	reg32 r1858 (rst, clk, r1857_out, r1858_out);
	reg32 r1859 (rst, clk, r1858_out, r1859_out);
	reg32 r1860 (rst, clk, r1859_out, r1860_out);
	reg32 r1861 (rst, clk, r1860_out, r1861_out);
	reg32 r1862 (rst, clk, r1861_out, r1862_out);
	reg32 r1863 (rst, clk, r1862_out, r1863_out);
	reg32 r1864 (rst, clk, r1863_out, r1864_out);
	reg32 r1865 (rst, clk, r1864_out, r1865_out);
	reg32 r1866 (rst, clk, r1865_out, r1866_out);
	reg32 r1867 (rst, clk, r1866_out, r1867_out);
	reg32 r1868 (rst, clk, r1867_out, r1868_out);
	reg32 r1869 (rst, clk, r1868_out, r1869_out);
	reg32 r1870 (rst, clk, r1869_out, r1870_out);
	reg32 r1871 (rst, clk, r1870_out, r1871_out);
	reg32 r1872 (rst, clk, r1871_out, r1872_out);
	reg32 r1873 (rst, clk, r1872_out, r1873_out);
	reg32 r1874 (rst, clk, r1873_out, r1874_out);
	reg32 r1875 (rst, clk, r1874_out, r1875_out);
	reg32 r1876 (rst, clk, r1875_out, r1876_out);
	reg32 r1877 (rst, clk, r1876_out, r1877_out);
	reg32 r1878 (rst, clk, r1877_out, r1878_out);
	reg32 r1879 (rst, clk, r1878_out, r1879_out);
	reg32 r1880 (rst, clk, r1879_out, r1880_out);
	reg32 r1881 (rst, clk, r1880_out, r1881_out);
	reg32 r1882 (rst, clk, r1881_out, r1882_out);
	reg32 r1883 (rst, clk, r1882_out, r1883_out);
	reg32 r1884 (rst, clk, r1883_out, r1884_out);
	reg32 r1885 (rst, clk, r1884_out, r1885_out);
	reg32 r1886 (rst, clk, r1885_out, r1886_out);
	reg32 r1887 (rst, clk, r1886_out, r1887_out);
	reg32 r1888 (rst, clk, r1887_out, r1888_out);
	reg32 r1889 (rst, clk, r1888_out, r1889_out);
	reg32 r1890 (rst, clk, r1889_out, r1890_out);
	reg32 r1891 (rst, clk, r1890_out, r1891_out);
	reg32 r1892 (rst, clk, r1891_out, r1892_out);
	reg32 r1893 (rst, clk, r1892_out, r1893_out);
	reg32 r1894 (rst, clk, r1893_out, r1894_out);
	reg32 r1895 (rst, clk, r1894_out, r1895_out);
	reg32 r1896 (rst, clk, r1895_out, r1896_out);
	reg32 r1897 (rst, clk, r1896_out, r1897_out);
	reg32 r1898 (rst, clk, r1897_out, r1898_out);
	reg32 r1899 (rst, clk, r1898_out, r1899_out);
	reg32 r1900 (rst, clk, r1899_out, r1900_out);
	reg32 r1901 (rst, clk, r1900_out, r1901_out);
	reg32 r1902 (rst, clk, r1901_out, r1902_out);
	reg32 r1903 (rst, clk, r1902_out, r1903_out);
	reg32 r1904 (rst, clk, r1903_out, r1904_out);
	reg32 r1905 (rst, clk, r1904_out, r1905_out);
	reg32 r1906 (rst, clk, r1905_out, r1906_out);
	reg32 r1907 (rst, clk, r1906_out, r1907_out);
	reg32 r1908 (rst, clk, r1907_out, r1908_out);
	reg32 r1909 (rst, clk, r1908_out, r1909_out);
	reg32 r1910 (rst, clk, r1909_out, r1910_out);
	reg32 r1911 (rst, clk, r1910_out, r1911_out);
	reg32 r1912 (rst, clk, r1911_out, r1912_out);
	reg32 r1913 (rst, clk, r1912_out, r1913_out);
	reg32 r1914 (rst, clk, r1913_out, r1914_out);
	reg32 r1915 (rst, clk, r1914_out, r1915_out);
	reg32 r1916 (rst, clk, r1915_out, r1916_out);
	reg32 r1917 (rst, clk, r1916_out, r1917_out);
	reg32 r1918 (rst, clk, r1917_out, r1918_out);
	reg32 r1919 (rst, clk, r1918_out, r1919_out);
	reg32 r1920 (rst, clk, r1919_out, r1920_out);
	reg32 r1921 (rst, clk, r1920_out, r1921_out);
	reg32 r1922 (rst, clk, r1921_out, r1922_out);
	reg32 r1923 (rst, clk, r1922_out, r1923_out);
	reg32 r1924 (rst, clk, r1923_out, r1924_out);
	reg32 r1925 (rst, clk, r1924_out, r1925_out);
	reg32 r1926 (rst, clk, r1925_out, r1926_out);
	reg32 r1927 (rst, clk, r1926_out, r1927_out);
	reg32 r1928 (rst, clk, r1927_out, r1928_out);
	reg32 r1929 (rst, clk, r1928_out, r1929_out);
	reg32 r1930 (rst, clk, r1929_out, r1930_out);
	reg32 r1931 (rst, clk, r1930_out, r1931_out);
	reg32 r1932 (rst, clk, r1931_out, r1932_out);
	reg32 r1933 (rst, clk, r1932_out, r1933_out);
	reg32 r1934 (rst, clk, r1933_out, r1934_out);
	reg32 r1935 (rst, clk, r1934_out, r1935_out);
	reg32 r1936 (rst, clk, r1935_out, r1936_out);
	reg32 r1937 (rst, clk, r1936_out, r1937_out);
	reg32 r1938 (rst, clk, r1937_out, r1938_out);
	reg32 r1939 (rst, clk, r1938_out, r1939_out);
	reg32 r1940 (rst, clk, r1939_out, r1940_out);
	reg32 r1941 (rst, clk, r1940_out, r1941_out);
	reg32 r1942 (rst, clk, r1941_out, r1942_out);
	reg32 r1943 (rst, clk, r1942_out, r1943_out);
	reg32 r1944 (rst, clk, r1943_out, r1944_out);
	reg32 r1945 (rst, clk, r1944_out, r1945_out);
	reg32 r1946 (rst, clk, r1945_out, r1946_out);
	reg32 r1947 (rst, clk, r1946_out, r1947_out);
	reg32 r1948 (rst, clk, r1947_out, r1948_out);
	reg32 r1949 (rst, clk, r1948_out, r1949_out);
	reg32 r1950 (rst, clk, r1949_out, r1950_out);
	reg32 r1951 (rst, clk, r1950_out, r1951_out);
	reg32 r1952 (rst, clk, r1951_out, r1952_out);
	reg32 r1953 (rst, clk, r1952_out, r1953_out);
	reg32 r1954 (rst, clk, r1953_out, r1954_out);
	reg32 r1955 (rst, clk, r1954_out, r1955_out);
	reg32 r1956 (rst, clk, r1955_out, r1956_out);
	reg32 r1957 (rst, clk, r1956_out, r1957_out);
	reg32 r1958 (rst, clk, r1957_out, r1958_out);
	reg32 r1959 (rst, clk, r1958_out, r1959_out);
	reg32 r1960 (rst, clk, r1959_out, r1960_out);
	reg32 r1961 (rst, clk, r1960_out, r1961_out);
	reg32 r1962 (rst, clk, r1961_out, r1962_out);
	reg32 r1963 (rst, clk, r1962_out, r1963_out);
	reg32 r1964 (rst, clk, r1963_out, r1964_out);
	reg32 r1965 (rst, clk, r1964_out, r1965_out);
	reg32 r1966 (rst, clk, r1965_out, r1966_out);
	reg32 r1967 (rst, clk, r1966_out, r1967_out);
	reg32 r1968 (rst, clk, r1967_out, r1968_out);
	reg32 r1969 (rst, clk, r1968_out, r1969_out);
	reg32 r1970 (rst, clk, r1969_out, r1970_out);
	reg32 r1971 (rst, clk, r1970_out, r1971_out);
	reg32 r1972 (rst, clk, r1971_out, r1972_out);
	reg32 r1973 (rst, clk, r1972_out, r1973_out);
	reg32 r1974 (rst, clk, r1973_out, r1974_out);
	reg32 r1975 (rst, clk, r1974_out, r1975_out);
	reg32 r1976 (rst, clk, r1975_out, r1976_out);
	reg32 r1977 (rst, clk, r1976_out, r1977_out);
	reg32 r1978 (rst, clk, r1977_out, r1978_out);
	reg32 r1979 (rst, clk, r1978_out, r1979_out);
	reg32 r1980 (rst, clk, r1979_out, r1980_out);
	reg32 r1981 (rst, clk, r1980_out, r1981_out);
	reg32 r1982 (rst, clk, r1981_out, r1982_out);
	reg32 r1983 (rst, clk, r1982_out, r1983_out);
	reg32 r1984 (rst, clk, r1983_out, r1984_out);
	reg32 r1985 (rst, clk, r1984_out, r1985_out);
	reg32 r1986 (rst, clk, r1985_out, r1986_out);
	reg32 r1987 (rst, clk, r1986_out, r1987_out);
	reg32 r1988 (rst, clk, r1987_out, r1988_out);
	reg32 r1989 (rst, clk, r1988_out, r1989_out);
	reg32 r1990 (rst, clk, r1989_out, r1990_out);
	reg32 r1991 (rst, clk, r1990_out, r1991_out);
	reg32 r1992 (rst, clk, r1991_out, r1992_out);
	reg32 r1993 (rst, clk, r1992_out, r1993_out);
	reg32 r1994 (rst, clk, r1993_out, r1994_out);
	reg32 r1995 (rst, clk, r1994_out, r1995_out);
	reg32 r1996 (rst, clk, r1995_out, r1996_out);
	reg32 r1997 (rst, clk, r1996_out, r1997_out);
	reg32 r1998 (rst, clk, r1997_out, r1998_out);
	reg32 r1999 (rst, clk, r1998_out, r1999_out);
	reg32 r2000 (rst, clk, r1999_out, r2000_out);
	reg32 r2001 (rst, clk, r2000_out, r2001_out);
	reg32 r2002 (rst, clk, r2001_out, r2002_out);
	reg32 r2003 (rst, clk, r2002_out, r2003_out);
	reg32 r2004 (rst, clk, r2003_out, r2004_out);
	reg32 r2005 (rst, clk, r2004_out, r2005_out);
	reg32 r2006 (rst, clk, r2005_out, r2006_out);
	reg32 r2007 (rst, clk, r2006_out, r2007_out);
	reg32 r2008 (rst, clk, r2007_out, r2008_out);
	reg32 r2009 (rst, clk, r2008_out, r2009_out);
	reg32 r2010 (rst, clk, r2009_out, r2010_out);
	reg32 r2011 (rst, clk, r2010_out, r2011_out);
	reg32 r2012 (rst, clk, r2011_out, r2012_out);
	reg32 r2013 (rst, clk, r2012_out, r2013_out);
	reg32 r2014 (rst, clk, r2013_out, r2014_out);
	reg32 r2015 (rst, clk, r2014_out, r2015_out);
	reg32 r2016 (rst, clk, r2015_out, r2016_out);
	reg32 r2017 (rst, clk, r2016_out, r2017_out);
	reg32 r2018 (rst, clk, r2017_out, r2018_out);
	reg32 r2019 (rst, clk, r2018_out, r2019_out);
	reg32 r2020 (rst, clk, r2019_out, r2020_out);
	reg32 r2021 (rst, clk, r2020_out, r2021_out);
	reg32 r2022 (rst, clk, r2021_out, r2022_out);
	reg32 r2023 (rst, clk, r2022_out, r2023_out);
	reg32 r2024 (rst, clk, r2023_out, r2024_out);
	reg32 r2025 (rst, clk, r2024_out, r2025_out);
	reg32 r2026 (rst, clk, r2025_out, r2026_out);
	reg32 r2027 (rst, clk, r2026_out, r2027_out);
	reg32 r2028 (rst, clk, r2027_out, r2028_out);
	reg32 r2029 (rst, clk, r2028_out, r2029_out);
	reg32 r2030 (rst, clk, r2029_out, r2030_out);
	reg32 r2031 (rst, clk, r2030_out, r2031_out);
	reg32 r2032 (rst, clk, r2031_out, r2032_out);
	reg32 r2033 (rst, clk, r2032_out, r2033_out);
	reg32 r2034 (rst, clk, r2033_out, r2034_out);
	reg32 r2035 (rst, clk, r2034_out, r2035_out);
	reg32 r2036 (rst, clk, r2035_out, r2036_out);
	reg32 r2037 (rst, clk, r2036_out, r2037_out);
	reg32 r2038 (rst, clk, r2037_out, r2038_out);
	reg32 r2039 (rst, clk, r2038_out, r2039_out);
	reg32 r2040 (rst, clk, r2039_out, r2040_out);
	reg32 r2041 (rst, clk, r2040_out, r2041_out);
	reg32 r2042 (rst, clk, r2041_out, r2042_out);
	reg32 r2043 (rst, clk, r2042_out, r2043_out);
	reg32 r2044 (rst, clk, r2043_out, r2044_out);
	reg32 r2045 (rst, clk, r2044_out, r2045_out);
	reg32 r2046 (rst, clk, r2045_out, r2046_out);
	reg32 r2047 (rst, clk, r2046_out, r2047_out);
	reg32 r2048 (rst, clk, r2047_out, r2048_out);
	reg32 r2049 (rst, clk, r2048_out, r2049_out);
	reg32 r2050 (rst, clk, r2049_out, r2050_out);
	reg32 r2051 (rst, clk, r2050_out, r2051_out);
	reg32 r2052 (rst, clk, r2051_out, r2052_out);
	reg32 r2053 (rst, clk, r2052_out, r2053_out);
	reg32 r2054 (rst, clk, r2053_out, r2054_out);
	reg32 r2055 (rst, clk, r2054_out, r2055_out);
	reg32 r2056 (rst, clk, r2055_out, r2056_out);
	reg32 r2057 (rst, clk, r2056_out, r2057_out);
	reg32 r2058 (rst, clk, r2057_out, r2058_out);
	reg32 r2059 (rst, clk, r2058_out, r2059_out);
	reg32 r2060 (rst, clk, r2059_out, r2060_out);
	reg32 r2061 (rst, clk, r2060_out, r2061_out);
	reg32 r2062 (rst, clk, r2061_out, r2062_out);
	reg32 r2063 (rst, clk, r2062_out, r2063_out);
	reg32 r2064 (rst, clk, r2063_out, r2064_out);
	reg32 r2065 (rst, clk, r2064_out, r2065_out);
	reg32 r2066 (rst, clk, r2065_out, r2066_out);
	reg32 r2067 (rst, clk, r2066_out, r2067_out);
	reg32 r2068 (rst, clk, r2067_out, r2068_out);
	reg32 r2069 (rst, clk, r2068_out, r2069_out);
	reg32 r2070 (rst, clk, r2069_out, r2070_out);
	reg32 r2071 (rst, clk, r2070_out, r2071_out);
	reg32 r2072 (rst, clk, r2071_out, r2072_out);
	reg32 r2073 (rst, clk, r2072_out, r2073_out);
	reg32 r2074 (rst, clk, r2073_out, r2074_out);
	reg32 r2075 (rst, clk, r2074_out, r2075_out);
	reg32 r2076 (rst, clk, r2075_out, r2076_out);
	reg32 r2077 (rst, clk, r2076_out, r2077_out);
	reg32 r2078 (rst, clk, r2077_out, r2078_out);
	reg32 r2079 (rst, clk, r2078_out, r2079_out);
	reg32 r2080 (rst, clk, r2079_out, r2080_out);
	reg32 r2081 (rst, clk, r2080_out, r2081_out);
	reg32 r2082 (rst, clk, r2081_out, r2082_out);
	reg32 r2083 (rst, clk, r2082_out, r2083_out);
	reg32 r2084 (rst, clk, r2083_out, r2084_out);
	reg32 r2085 (rst, clk, r2084_out, r2085_out);
	reg32 r2086 (rst, clk, r2085_out, r2086_out);
	reg32 r2087 (rst, clk, r2086_out, r2087_out);
	reg32 r2088 (rst, clk, r2087_out, r2088_out);
	reg32 r2089 (rst, clk, r2088_out, r2089_out);
	reg32 r2090 (rst, clk, r2089_out, r2090_out);
	reg32 r2091 (rst, clk, r2090_out, r2091_out);
	reg32 r2092 (rst, clk, r2091_out, r2092_out);
	reg32 r2093 (rst, clk, r2092_out, r2093_out);
	reg32 r2094 (rst, clk, r2093_out, r2094_out);
	reg32 r2095 (rst, clk, r2094_out, r2095_out);
	reg32 r2096 (rst, clk, r2095_out, r2096_out);
	reg32 r2097 (rst, clk, r2096_out, r2097_out);
	reg32 r2098 (rst, clk, r2097_out, r2098_out);
	reg32 r2099 (rst, clk, r2098_out, r2099_out);
	reg32 r2100 (rst, clk, r2099_out, r2100_out);
	reg32 r2101 (rst, clk, r2100_out, r2101_out);
	reg32 r2102 (rst, clk, r2101_out, r2102_out);
	reg32 r2103 (rst, clk, r2102_out, r2103_out);
	reg32 r2104 (rst, clk, r2103_out, r2104_out);
	reg32 r2105 (rst, clk, r2104_out, r2105_out);
	reg32 r2106 (rst, clk, r2105_out, r2106_out);
	reg32 r2107 (rst, clk, r2106_out, r2107_out);
	reg32 r2108 (rst, clk, r2107_out, r2108_out);
	reg32 r2109 (rst, clk, r2108_out, r2109_out);
	reg32 r2110 (rst, clk, r2109_out, r2110_out);
	reg32 r2111 (rst, clk, r2110_out, r2111_out);
	reg32 r2112 (rst, clk, r2111_out, r2112_out);
	reg32 r2113 (rst, clk, r2112_out, r2113_out);
	reg32 r2114 (rst, clk, r2113_out, r2114_out);
	reg32 r2115 (rst, clk, r2114_out, r2115_out);
	reg32 r2116 (rst, clk, r2115_out, r2116_out);
	reg32 r2117 (rst, clk, r2116_out, r2117_out);
	reg32 r2118 (rst, clk, r2117_out, r2118_out);
	reg32 r2119 (rst, clk, r2118_out, r2119_out);
	reg32 r2120 (rst, clk, r2119_out, r2120_out);
	reg32 r2121 (rst, clk, r2120_out, r2121_out);
	reg32 r2122 (rst, clk, r2121_out, r2122_out);
	reg32 r2123 (rst, clk, r2122_out, r2123_out);
	reg32 r2124 (rst, clk, r2123_out, r2124_out);
	reg32 r2125 (rst, clk, r2124_out, r2125_out);
	reg32 r2126 (rst, clk, r2125_out, r2126_out);
	reg32 r2127 (rst, clk, r2126_out, r2127_out);
	reg32 r2128 (rst, clk, r2127_out, r2128_out);
	reg32 r2129 (rst, clk, r2128_out, r2129_out);
	reg32 r2130 (rst, clk, r2129_out, r2130_out);
	reg32 r2131 (rst, clk, r2130_out, r2131_out);
	reg32 r2132 (rst, clk, r2131_out, r2132_out);
	reg32 r2133 (rst, clk, r2132_out, r2133_out);
	reg32 r2134 (rst, clk, r2133_out, r2134_out);
	reg32 r2135 (rst, clk, r2134_out, r2135_out);
	reg32 r2136 (rst, clk, r2135_out, r2136_out);
	reg32 r2137 (rst, clk, r2136_out, r2137_out);
	reg32 r2138 (rst, clk, r2137_out, r2138_out);
	reg32 r2139 (rst, clk, r2138_out, r2139_out);
	reg32 r2140 (rst, clk, r2139_out, r2140_out);
	reg32 r2141 (rst, clk, r2140_out, r2141_out);
	reg32 r2142 (rst, clk, r2141_out, r2142_out);
	reg32 r2143 (rst, clk, r2142_out, r2143_out);
	reg32 r2144 (rst, clk, r2143_out, r2144_out);
	reg32 r2145 (rst, clk, r2144_out, r2145_out);
	reg32 r2146 (rst, clk, r2145_out, r2146_out);
	reg32 r2147 (rst, clk, r2146_out, r2147_out);
	reg32 r2148 (rst, clk, r2147_out, r2148_out);
	reg32 r2149 (rst, clk, r2148_out, r2149_out);
	reg32 r2150 (rst, clk, r2149_out, r2150_out);
	reg32 r2151 (rst, clk, r2150_out, r2151_out);
	reg32 r2152 (rst, clk, r2151_out, r2152_out);
	reg32 r2153 (rst, clk, r2152_out, r2153_out);
	reg32 r2154 (rst, clk, r2153_out, r2154_out);
	reg32 r2155 (rst, clk, r2154_out, r2155_out);
	reg32 r2156 (rst, clk, r2155_out, r2156_out);
	reg32 r2157 (rst, clk, r2156_out, r2157_out);
	reg32 r2158 (rst, clk, r2157_out, r2158_out);
	reg32 r2159 (rst, clk, r2158_out, r2159_out);
	reg32 r2160 (rst, clk, r2159_out, r2160_out);
	reg32 r2161 (rst, clk, r2160_out, r2161_out);
	reg32 r2162 (rst, clk, r2161_out, r2162_out);
	reg32 r2163 (rst, clk, r2162_out, r2163_out);
	reg32 r2164 (rst, clk, r2163_out, r2164_out);
	reg32 r2165 (rst, clk, r2164_out, r2165_out);
	reg32 r2166 (rst, clk, r2165_out, r2166_out);
	reg32 r2167 (rst, clk, r2166_out, r2167_out);
	reg32 r2168 (rst, clk, r2167_out, r2168_out);
	reg32 r2169 (rst, clk, r2168_out, r2169_out);
	reg32 r2170 (rst, clk, r2169_out, r2170_out);
	reg32 r2171 (rst, clk, r2170_out, r2171_out);
	reg32 r2172 (rst, clk, r2171_out, r2172_out);
	reg32 r2173 (rst, clk, r2172_out, r2173_out);
	reg32 r2174 (rst, clk, r2173_out, r2174_out);
	reg32 r2175 (rst, clk, r2174_out, r2175_out);
	reg32 r2176 (rst, clk, r2175_out, r2176_out);
	reg32 r2177 (rst, clk, r2176_out, r2177_out);
	reg32 r2178 (rst, clk, r2177_out, r2178_out);
	reg32 r2179 (rst, clk, r2178_out, r2179_out);
	reg32 r2180 (rst, clk, r2179_out, r2180_out);
	reg32 r2181 (rst, clk, r2180_out, r2181_out);
	reg32 r2182 (rst, clk, r2181_out, r2182_out);
	reg32 r2183 (rst, clk, r2182_out, r2183_out);
	reg32 r2184 (rst, clk, r2183_out, r2184_out);
	reg32 r2185 (rst, clk, r2184_out, r2185_out);
	reg32 r2186 (rst, clk, r2185_out, r2186_out);
	reg32 r2187 (rst, clk, r2186_out, r2187_out);
	reg32 r2188 (rst, clk, r2187_out, r2188_out);
	reg32 r2189 (rst, clk, r2188_out, r2189_out);
	reg32 r2190 (rst, clk, r2189_out, r2190_out);
	reg32 r2191 (rst, clk, r2190_out, r2191_out);
	reg32 r2192 (rst, clk, r2191_out, r2192_out);
	reg32 r2193 (rst, clk, r2192_out, r2193_out);
	reg32 r2194 (rst, clk, r2193_out, r2194_out);
	reg32 r2195 (rst, clk, r2194_out, r2195_out);
	reg32 r2196 (rst, clk, r2195_out, r2196_out);
	reg32 r2197 (rst, clk, r2196_out, r2197_out);
	reg32 r2198 (rst, clk, r2197_out, r2198_out);
	reg32 r2199 (rst, clk, r2198_out, r2199_out);
	reg32 r2200 (rst, clk, r2199_out, r2200_out);
	reg32 r2201 (rst, clk, r2200_out, r2201_out);
	reg32 r2202 (rst, clk, r2201_out, r2202_out);
	reg32 r2203 (rst, clk, r2202_out, r2203_out);
	reg32 r2204 (rst, clk, r2203_out, r2204_out);
	reg32 r2205 (rst, clk, r2204_out, r2205_out);
	reg32 r2206 (rst, clk, r2205_out, r2206_out);
	reg32 r2207 (rst, clk, r2206_out, r2207_out);
	reg32 r2208 (rst, clk, r2207_out, r2208_out);
	reg32 r2209 (rst, clk, r2208_out, r2209_out);
	reg32 r2210 (rst, clk, r2209_out, r2210_out);
	reg32 r2211 (rst, clk, r2210_out, r2211_out);
	reg32 r2212 (rst, clk, r2211_out, r2212_out);
	reg32 r2213 (rst, clk, r2212_out, r2213_out);
	reg32 r2214 (rst, clk, r2213_out, r2214_out);
	reg32 r2215 (rst, clk, r2214_out, r2215_out);
	reg32 r2216 (rst, clk, r2215_out, r2216_out);
	reg32 r2217 (rst, clk, r2216_out, r2217_out);
	reg32 r2218 (rst, clk, r2217_out, r2218_out);
	reg32 r2219 (rst, clk, r2218_out, r2219_out);
	reg32 r2220 (rst, clk, r2219_out, r2220_out);
	reg32 r2221 (rst, clk, r2220_out, r2221_out);
	reg32 r2222 (rst, clk, r2221_out, r2222_out);
	reg32 r2223 (rst, clk, r2222_out, r2223_out);
	reg32 r2224 (rst, clk, r2223_out, r2224_out);
	reg32 r2225 (rst, clk, r2224_out, r2225_out);
	reg32 r2226 (rst, clk, r2225_out, r2226_out);
	reg32 r2227 (rst, clk, r2226_out, r2227_out);
	reg32 r2228 (rst, clk, r2227_out, r2228_out);
	reg32 r2229 (rst, clk, r2228_out, r2229_out);
	reg32 r2230 (rst, clk, r2229_out, r2230_out);
	reg32 r2231 (rst, clk, r2230_out, r2231_out);
	reg32 r2232 (rst, clk, r2231_out, r2232_out);
	reg32 r2233 (rst, clk, r2232_out, r2233_out);
	reg32 r2234 (rst, clk, r2233_out, r2234_out);
	reg32 r2235 (rst, clk, r2234_out, r2235_out);
	reg32 r2236 (rst, clk, r2235_out, r2236_out);
	reg32 r2237 (rst, clk, r2236_out, r2237_out);
	reg32 r2238 (rst, clk, r2237_out, r2238_out);
	reg32 r2239 (rst, clk, r2238_out, r2239_out);
	reg32 r2240 (rst, clk, r2239_out, r2240_out);
	reg32 r2241 (rst, clk, r2240_out, r2241_out);
	reg32 r2242 (rst, clk, r2241_out, r2242_out);
	reg32 r2243 (rst, clk, r2242_out, r2243_out);
	reg32 r2244 (rst, clk, r2243_out, r2244_out);
	reg32 r2245 (rst, clk, r2244_out, r2245_out);
	reg32 r2246 (rst, clk, r2245_out, r2246_out);
	reg32 r2247 (rst, clk, r2246_out, r2247_out);
	reg32 r2248 (rst, clk, r2247_out, r2248_out);
	reg32 r2249 (rst, clk, r2248_out, r2249_out);
	reg32 r2250 (rst, clk, r2249_out, r2250_out);
	reg32 r2251 (rst, clk, r2250_out, r2251_out);
	reg32 r2252 (rst, clk, r2251_out, r2252_out);
	reg32 r2253 (rst, clk, r2252_out, r2253_out);
	reg32 r2254 (rst, clk, r2253_out, r2254_out);
	reg32 r2255 (rst, clk, r2254_out, r2255_out);
	reg32 r2256 (rst, clk, r2255_out, r2256_out);
	reg32 r2257 (rst, clk, r2256_out, r2257_out);
	reg32 r2258 (rst, clk, r2257_out, r2258_out);
	reg32 r2259 (rst, clk, r2258_out, r2259_out);
	reg32 r2260 (rst, clk, r2259_out, r2260_out);
	reg32 r2261 (rst, clk, r2260_out, r2261_out);
	reg32 r2262 (rst, clk, r2261_out, r2262_out);
	reg32 r2263 (rst, clk, r2262_out, r2263_out);
	reg32 r2264 (rst, clk, r2263_out, r2264_out);
	reg32 r2265 (rst, clk, r2264_out, r2265_out);
	reg32 r2266 (rst, clk, r2265_out, r2266_out);
	reg32 r2267 (rst, clk, r2266_out, r2267_out);
	reg32 r2268 (rst, clk, r2267_out, r2268_out);
	reg32 r2269 (rst, clk, r2268_out, r2269_out);
	reg32 r2270 (rst, clk, r2269_out, r2270_out);
	reg32 r2271 (rst, clk, r2270_out, r2271_out);
	reg32 r2272 (rst, clk, r2271_out, r2272_out);
	reg32 r2273 (rst, clk, r2272_out, r2273_out);
	reg32 r2274 (rst, clk, r2273_out, r2274_out);
	reg32 r2275 (rst, clk, r2274_out, r2275_out);
	reg32 r2276 (rst, clk, r2275_out, r2276_out);
	reg32 r2277 (rst, clk, r2276_out, r2277_out);
	reg32 r2278 (rst, clk, r2277_out, r2278_out);
	reg32 r2279 (rst, clk, r2278_out, r2279_out);
	reg32 r2280 (rst, clk, r2279_out, r2280_out);
	reg32 r2281 (rst, clk, r2280_out, r2281_out);
	reg32 r2282 (rst, clk, r2281_out, r2282_out);
	reg32 r2283 (rst, clk, r2282_out, r2283_out);
	reg32 r2284 (rst, clk, r2283_out, r2284_out);
	reg32 r2285 (rst, clk, r2284_out, r2285_out);
	reg32 r2286 (rst, clk, r2285_out, r2286_out);
	reg32 r2287 (rst, clk, r2286_out, r2287_out);
	reg32 r2288 (rst, clk, r2287_out, r2288_out);
	reg32 r2289 (rst, clk, r2288_out, r2289_out);
	reg32 r2290 (rst, clk, r2289_out, r2290_out);
	reg32 r2291 (rst, clk, r2290_out, r2291_out);
	reg32 r2292 (rst, clk, r2291_out, r2292_out);
	reg32 r2293 (rst, clk, r2292_out, r2293_out);
	reg32 r2294 (rst, clk, r2293_out, r2294_out);
	reg32 r2295 (rst, clk, r2294_out, r2295_out);
	reg32 r2296 (rst, clk, r2295_out, r2296_out);
	reg32 r2297 (rst, clk, r2296_out, r2297_out);
	reg32 r2298 (rst, clk, r2297_out, r2298_out);
	reg32 r2299 (rst, clk, r2298_out, r2299_out);
	reg32 r2300 (rst, clk, r2299_out, r2300_out);
	reg32 r2301 (rst, clk, r2300_out, r2301_out);
	reg32 r2302 (rst, clk, r2301_out, r2302_out);
	reg32 r2303 (rst, clk, r2302_out, r2303_out);
	reg32 r2304 (rst, clk, r2303_out, r2304_out);
	reg32 r2305 (rst, clk, r2304_out, r2305_out);
	reg32 r2306 (rst, clk, r2305_out, r2306_out);
	reg32 r2307 (rst, clk, r2306_out, r2307_out);
	reg32 r2308 (rst, clk, r2307_out, r2308_out);
	reg32 r2309 (rst, clk, r2308_out, r2309_out);
	reg32 r2310 (rst, clk, r2309_out, r2310_out);
	reg32 r2311 (rst, clk, r2310_out, r2311_out);
	reg32 r2312 (rst, clk, r2311_out, r2312_out);
	reg32 r2313 (rst, clk, r2312_out, r2313_out);
	reg32 r2314 (rst, clk, r2313_out, r2314_out);
	reg32 r2315 (rst, clk, r2314_out, r2315_out);
	reg32 r2316 (rst, clk, r2315_out, r2316_out);
	reg32 r2317 (rst, clk, r2316_out, r2317_out);
	reg32 r2318 (rst, clk, r2317_out, r2318_out);
	reg32 r2319 (rst, clk, r2318_out, r2319_out);
	reg32 r2320 (rst, clk, r2319_out, r2320_out);
	reg32 r2321 (rst, clk, r2320_out, r2321_out);
	reg32 r2322 (rst, clk, r2321_out, r2322_out);
	reg32 r2323 (rst, clk, r2322_out, r2323_out);
	reg32 r2324 (rst, clk, r2323_out, r2324_out);
	reg32 r2325 (rst, clk, r2324_out, r2325_out);
	reg32 r2326 (rst, clk, r2325_out, r2326_out);
	reg32 r2327 (rst, clk, r2326_out, r2327_out);
	reg32 r2328 (rst, clk, r2327_out, r2328_out);
	reg32 r2329 (rst, clk, r2328_out, r2329_out);
	reg32 r2330 (rst, clk, r2329_out, r2330_out);
	reg32 r2331 (rst, clk, r2330_out, r2331_out);
	reg32 r2332 (rst, clk, r2331_out, r2332_out);
	reg32 r2333 (rst, clk, r2332_out, r2333_out);
	reg32 r2334 (rst, clk, r2333_out, r2334_out);
	reg32 r2335 (rst, clk, r2334_out, r2335_out);
	reg32 r2336 (rst, clk, r2335_out, r2336_out);
	reg32 r2337 (rst, clk, r2336_out, r2337_out);
	reg32 r2338 (rst, clk, r2337_out, r2338_out);
	reg32 r2339 (rst, clk, r2338_out, r2339_out);
	reg32 r2340 (rst, clk, r2339_out, r2340_out);
	reg32 r2341 (rst, clk, r2340_out, r2341_out);
	reg32 r2342 (rst, clk, r2341_out, r2342_out);
	reg32 r2343 (rst, clk, r2342_out, r2343_out);
	reg32 r2344 (rst, clk, r2343_out, r2344_out);
	reg32 r2345 (rst, clk, r2344_out, r2345_out);
	reg32 r2346 (rst, clk, r2345_out, r2346_out);
	reg32 r2347 (rst, clk, r2346_out, r2347_out);
	reg32 r2348 (rst, clk, r2347_out, r2348_out);
	reg32 r2349 (rst, clk, r2348_out, r2349_out);
	reg32 r2350 (rst, clk, r2349_out, r2350_out);
	reg32 r2351 (rst, clk, r2350_out, r2351_out);
	reg32 r2352 (rst, clk, r2351_out, r2352_out);
	reg32 r2353 (rst, clk, r2352_out, r2353_out);
	reg32 r2354 (rst, clk, r2353_out, r2354_out);
	reg32 r2355 (rst, clk, r2354_out, r2355_out);
	reg32 r2356 (rst, clk, r2355_out, r2356_out);
	reg32 r2357 (rst, clk, r2356_out, r2357_out);
	reg32 r2358 (rst, clk, r2357_out, r2358_out);
	reg32 r2359 (rst, clk, r2358_out, r2359_out);
	reg32 r2360 (rst, clk, r2359_out, r2360_out);
	reg32 r2361 (rst, clk, r2360_out, r2361_out);
	reg32 r2362 (rst, clk, r2361_out, r2362_out);
	reg32 r2363 (rst, clk, r2362_out, r2363_out);
	reg32 r2364 (rst, clk, r2363_out, r2364_out);
	reg32 r2365 (rst, clk, r2364_out, r2365_out);
	reg32 r2366 (rst, clk, r2365_out, r2366_out);
	reg32 r2367 (rst, clk, r2366_out, r2367_out);
	reg32 r2368 (rst, clk, r2367_out, r2368_out);
	reg32 r2369 (rst, clk, r2368_out, r2369_out);
	reg32 r2370 (rst, clk, r2369_out, r2370_out);
	reg32 r2371 (rst, clk, r2370_out, r2371_out);
	reg32 r2372 (rst, clk, r2371_out, r2372_out);
	reg32 r2373 (rst, clk, r2372_out, r2373_out);
	reg32 r2374 (rst, clk, r2373_out, r2374_out);
	reg32 r2375 (rst, clk, r2374_out, r2375_out);
	reg32 r2376 (rst, clk, r2375_out, r2376_out);
	reg32 r2377 (rst, clk, r2376_out, r2377_out);
	reg32 r2378 (rst, clk, r2377_out, r2378_out);
	reg32 r2379 (rst, clk, r2378_out, r2379_out);
	reg32 r2380 (rst, clk, r2379_out, r2380_out);
	reg32 r2381 (rst, clk, r2380_out, r2381_out);
	reg32 r2382 (rst, clk, r2381_out, r2382_out);
	reg32 r2383 (rst, clk, r2382_out, r2383_out);
	reg32 r2384 (rst, clk, r2383_out, r2384_out);
	reg32 r2385 (rst, clk, r2384_out, r2385_out);
	reg32 r2386 (rst, clk, r2385_out, r2386_out);
	reg32 r2387 (rst, clk, r2386_out, r2387_out);
	reg32 r2388 (rst, clk, r2387_out, r2388_out);
	reg32 r2389 (rst, clk, r2388_out, r2389_out);
	reg32 r2390 (rst, clk, r2389_out, r2390_out);
	reg32 r2391 (rst, clk, r2390_out, r2391_out);
	reg32 r2392 (rst, clk, r2391_out, r2392_out);
	reg32 r2393 (rst, clk, r2392_out, r2393_out);
	reg32 r2394 (rst, clk, r2393_out, r2394_out);
	reg32 r2395 (rst, clk, r2394_out, r2395_out);
	reg32 r2396 (rst, clk, r2395_out, r2396_out);
	reg32 r2397 (rst, clk, r2396_out, r2397_out);
	reg32 r2398 (rst, clk, r2397_out, r2398_out);
	reg32 r2399 (rst, clk, r2398_out, r2399_out);
	reg32 r2400 (rst, clk, r2399_out, r2400_out);
	reg32 r2401 (rst, clk, r2400_out, r2401_out);
	reg32 r2402 (rst, clk, r2401_out, r2402_out);
	reg32 r2403 (rst, clk, r2402_out, r2403_out);
	reg32 r2404 (rst, clk, r2403_out, r2404_out);
	reg32 r2405 (rst, clk, r2404_out, r2405_out);
	reg32 r2406 (rst, clk, r2405_out, r2406_out);
	reg32 r2407 (rst, clk, r2406_out, r2407_out);
	reg32 r2408 (rst, clk, r2407_out, r2408_out);
	reg32 r2409 (rst, clk, r2408_out, r2409_out);
	reg32 r2410 (rst, clk, r2409_out, r2410_out);
	reg32 r2411 (rst, clk, r2410_out, r2411_out);
	reg32 r2412 (rst, clk, r2411_out, r2412_out);
	reg32 r2413 (rst, clk, r2412_out, r2413_out);
	reg32 r2414 (rst, clk, r2413_out, r2414_out);
	reg32 r2415 (rst, clk, r2414_out, r2415_out);
	reg32 r2416 (rst, clk, r2415_out, r2416_out);
	reg32 r2417 (rst, clk, r2416_out, r2417_out);
	reg32 r2418 (rst, clk, r2417_out, r2418_out);
	reg32 r2419 (rst, clk, r2418_out, r2419_out);
	reg32 r2420 (rst, clk, r2419_out, r2420_out);
	reg32 r2421 (rst, clk, r2420_out, r2421_out);
	reg32 r2422 (rst, clk, r2421_out, r2422_out);
	reg32 r2423 (rst, clk, r2422_out, r2423_out);
	reg32 r2424 (rst, clk, r2423_out, r2424_out);
	reg32 r2425 (rst, clk, r2424_out, r2425_out);
	reg32 r2426 (rst, clk, r2425_out, r2426_out);
	reg32 r2427 (rst, clk, r2426_out, r2427_out);
	reg32 r2428 (rst, clk, r2427_out, r2428_out);
	reg32 r2429 (rst, clk, r2428_out, r2429_out);
	reg32 r2430 (rst, clk, r2429_out, r2430_out);
	reg32 r2431 (rst, clk, r2430_out, r2431_out);
	reg32 r2432 (rst, clk, r2431_out, r2432_out);
	reg32 r2433 (rst, clk, r2432_out, r2433_out);
	reg32 r2434 (rst, clk, r2433_out, r2434_out);
	reg32 r2435 (rst, clk, r2434_out, r2435_out);
	reg32 r2436 (rst, clk, r2435_out, r2436_out);
	reg32 r2437 (rst, clk, r2436_out, r2437_out);
	reg32 r2438 (rst, clk, r2437_out, r2438_out);
	reg32 r2439 (rst, clk, r2438_out, r2439_out);
	reg32 r2440 (rst, clk, r2439_out, r2440_out);
	reg32 r2441 (rst, clk, r2440_out, r2441_out);
	reg32 r2442 (rst, clk, r2441_out, r2442_out);
	reg32 r2443 (rst, clk, r2442_out, r2443_out);
	reg32 r2444 (rst, clk, r2443_out, r2444_out);
	reg32 r2445 (rst, clk, r2444_out, r2445_out);
	reg32 r2446 (rst, clk, r2445_out, r2446_out);
	reg32 r2447 (rst, clk, r2446_out, r2447_out);
	reg32 r2448 (rst, clk, r2447_out, r2448_out);
	reg32 r2449 (rst, clk, r2448_out, r2449_out);
	reg32 r2450 (rst, clk, r2449_out, r2450_out);
	reg32 r2451 (rst, clk, r2450_out, r2451_out);
	reg32 r2452 (rst, clk, r2451_out, r2452_out);
	reg32 r2453 (rst, clk, r2452_out, r2453_out);
	reg32 r2454 (rst, clk, r2453_out, r2454_out);
	reg32 r2455 (rst, clk, r2454_out, r2455_out);
	reg32 r2456 (rst, clk, r2455_out, r2456_out);
	reg32 r2457 (rst, clk, r2456_out, r2457_out);
	reg32 r2458 (rst, clk, r2457_out, r2458_out);
	reg32 r2459 (rst, clk, r2458_out, r2459_out);
	reg32 r2460 (rst, clk, r2459_out, r2460_out);
	reg32 r2461 (rst, clk, r2460_out, r2461_out);
	reg32 r2462 (rst, clk, r2461_out, r2462_out);
	reg32 r2463 (rst, clk, r2462_out, r2463_out);
	reg32 r2464 (rst, clk, r2463_out, r2464_out);
	reg32 r2465 (rst, clk, r2464_out, r2465_out);
	reg32 r2466 (rst, clk, r2465_out, r2466_out);
	reg32 r2467 (rst, clk, r2466_out, r2467_out);
	reg32 r2468 (rst, clk, r2467_out, r2468_out);
	reg32 r2469 (rst, clk, r2468_out, r2469_out);
	reg32 r2470 (rst, clk, r2469_out, r2470_out);
	reg32 r2471 (rst, clk, r2470_out, r2471_out);
	reg32 r2472 (rst, clk, r2471_out, r2472_out);
	reg32 r2473 (rst, clk, r2472_out, r2473_out);
	reg32 r2474 (rst, clk, r2473_out, r2474_out);
	reg32 r2475 (rst, clk, r2474_out, r2475_out);
	reg32 r2476 (rst, clk, r2475_out, r2476_out);
	reg32 r2477 (rst, clk, r2476_out, r2477_out);
	reg32 r2478 (rst, clk, r2477_out, r2478_out);
	reg32 r2479 (rst, clk, r2478_out, r2479_out);
	reg32 r2480 (rst, clk, r2479_out, r2480_out);
	reg32 r2481 (rst, clk, r2480_out, r2481_out);
	reg32 r2482 (rst, clk, r2481_out, r2482_out);
	reg32 r2483 (rst, clk, r2482_out, r2483_out);
	reg32 r2484 (rst, clk, r2483_out, r2484_out);
	reg32 r2485 (rst, clk, r2484_out, r2485_out);
	reg32 r2486 (rst, clk, r2485_out, r2486_out);
	reg32 r2487 (rst, clk, r2486_out, r2487_out);
	reg32 r2488 (rst, clk, r2487_out, r2488_out);
	reg32 r2489 (rst, clk, r2488_out, r2489_out);
	reg32 r2490 (rst, clk, r2489_out, r2490_out);
	reg32 r2491 (rst, clk, r2490_out, r2491_out);
	reg32 r2492 (rst, clk, r2491_out, r2492_out);
	reg32 r2493 (rst, clk, r2492_out, r2493_out);
	reg32 r2494 (rst, clk, r2493_out, r2494_out);
	reg32 r2495 (rst, clk, r2494_out, r2495_out);
	reg32 r2496 (rst, clk, r2495_out, r2496_out);
	reg32 r2497 (rst, clk, r2496_out, r2497_out);
	reg32 r2498 (rst, clk, r2497_out, r2498_out);
	reg32 r2499 (rst, clk, r2498_out, r2499_out);
	reg32 r2500 (rst, clk, r2499_out, r2500_out);
	reg32 r2501 (rst, clk, r2500_out, r2501_out);
	reg32 r2502 (rst, clk, r2501_out, r2502_out);
	reg32 r2503 (rst, clk, r2502_out, r2503_out);
	reg32 r2504 (rst, clk, r2503_out, r2504_out);
	reg32 r2505 (rst, clk, r2504_out, r2505_out);
	reg32 r2506 (rst, clk, r2505_out, r2506_out);
	reg32 r2507 (rst, clk, r2506_out, r2507_out);
	reg32 r2508 (rst, clk, r2507_out, r2508_out);
	reg32 r2509 (rst, clk, r2508_out, r2509_out);
	reg32 r2510 (rst, clk, r2509_out, r2510_out);
	reg32 r2511 (rst, clk, r2510_out, r2511_out);
	reg32 r2512 (rst, clk, r2511_out, r2512_out);
	reg32 r2513 (rst, clk, r2512_out, r2513_out);
	reg32 r2514 (rst, clk, r2513_out, r2514_out);
	reg32 r2515 (rst, clk, r2514_out, r2515_out);
	reg32 r2516 (rst, clk, r2515_out, r2516_out);
	reg32 r2517 (rst, clk, r2516_out, r2517_out);
	reg32 r2518 (rst, clk, r2517_out, r2518_out);
	reg32 r2519 (rst, clk, r2518_out, r2519_out);
	reg32 r2520 (rst, clk, r2519_out, r2520_out);
	reg32 r2521 (rst, clk, r2520_out, r2521_out);
	reg32 r2522 (rst, clk, r2521_out, r2522_out);
	reg32 r2523 (rst, clk, r2522_out, r2523_out);
	reg32 r2524 (rst, clk, r2523_out, r2524_out);
	reg32 r2525 (rst, clk, r2524_out, r2525_out);
	reg32 r2526 (rst, clk, r2525_out, r2526_out);
	reg32 r2527 (rst, clk, r2526_out, r2527_out);
	reg32 r2528 (rst, clk, r2527_out, r2528_out);
	reg32 r2529 (rst, clk, r2528_out, r2529_out);
	reg32 r2530 (rst, clk, r2529_out, r2530_out);
	reg32 r2531 (rst, clk, r2530_out, r2531_out);
	reg32 r2532 (rst, clk, r2531_out, r2532_out);
	reg32 r2533 (rst, clk, r2532_out, r2533_out);
	reg32 r2534 (rst, clk, r2533_out, r2534_out);
	reg32 r2535 (rst, clk, r2534_out, r2535_out);
	reg32 r2536 (rst, clk, r2535_out, r2536_out);
	reg32 r2537 (rst, clk, r2536_out, r2537_out);
	reg32 r2538 (rst, clk, r2537_out, r2538_out);
	reg32 r2539 (rst, clk, r2538_out, r2539_out);
	reg32 r2540 (rst, clk, r2539_out, r2540_out);
	reg32 r2541 (rst, clk, r2540_out, r2541_out);
	reg32 r2542 (rst, clk, r2541_out, r2542_out);
	reg32 r2543 (rst, clk, r2542_out, r2543_out);
	reg32 r2544 (rst, clk, r2543_out, r2544_out);
	reg32 r2545 (rst, clk, r2544_out, r2545_out);
	reg32 r2546 (rst, clk, r2545_out, r2546_out);
	reg32 r2547 (rst, clk, r2546_out, r2547_out);
	reg32 r2548 (rst, clk, r2547_out, r2548_out);
	reg32 r2549 (rst, clk, r2548_out, r2549_out);
	reg32 r2550 (rst, clk, r2549_out, r2550_out);
	reg32 r2551 (rst, clk, r2550_out, r2551_out);
	reg32 r2552 (rst, clk, r2551_out, r2552_out);
	reg32 r2553 (rst, clk, r2552_out, r2553_out);
	reg32 r2554 (rst, clk, r2553_out, r2554_out);
	reg32 r2555 (rst, clk, r2554_out, r2555_out);
	reg32 r2556 (rst, clk, r2555_out, r2556_out);
	reg32 r2557 (rst, clk, r2556_out, r2557_out);
	reg32 r2558 (rst, clk, r2557_out, r2558_out);
	reg32 r2559 (rst, clk, r2558_out, r2559_out);
	reg32 r2560 (rst, clk, r2559_out, r2560_out);
	reg32 r2561 (rst, clk, r2560_out, r2561_out);
	reg32 r2562 (rst, clk, r2561_out, r2562_out);
	reg32 r2563 (rst, clk, r2562_out, r2563_out);
	reg32 r2564 (rst, clk, r2563_out, r2564_out);
	reg32 r2565 (rst, clk, r2564_out, r2565_out);
	reg32 r2566 (rst, clk, r2565_out, r2566_out);
	reg32 r2567 (rst, clk, r2566_out, r2567_out);
	reg32 r2568 (rst, clk, r2567_out, r2568_out);
	reg32 r2569 (rst, clk, r2568_out, r2569_out);
	reg32 r2570 (rst, clk, r2569_out, r2570_out);
	reg32 r2571 (rst, clk, r2570_out, r2571_out);
	reg32 r2572 (rst, clk, r2571_out, r2572_out);
	reg32 r2573 (rst, clk, r2572_out, r2573_out);
	reg32 r2574 (rst, clk, r2573_out, r2574_out);
	reg32 r2575 (rst, clk, r2574_out, r2575_out);
	reg32 r2576 (rst, clk, r2575_out, r2576_out);
	reg32 r2577 (rst, clk, r2576_out, r2577_out);
	reg32 r2578 (rst, clk, r2577_out, r2578_out);
	reg32 r2579 (rst, clk, r2578_out, r2579_out);
	reg32 r2580 (rst, clk, r2579_out, r2580_out);
	reg32 r2581 (rst, clk, r2580_out, r2581_out);
	reg32 r2582 (rst, clk, r2581_out, r2582_out);
	reg32 r2583 (rst, clk, r2582_out, r2583_out);
	reg32 r2584 (rst, clk, r2583_out, r2584_out);
	reg32 r2585 (rst, clk, r2584_out, r2585_out);
	reg32 r2586 (rst, clk, r2585_out, r2586_out);
	reg32 r2587 (rst, clk, r2586_out, r2587_out);
	reg32 r2588 (rst, clk, r2587_out, r2588_out);
	reg32 r2589 (rst, clk, r2588_out, r2589_out);
	reg32 r2590 (rst, clk, r2589_out, r2590_out);
	reg32 r2591 (rst, clk, r2590_out, r2591_out);
	reg32 r2592 (rst, clk, r2591_out, r2592_out);
	reg32 r2593 (rst, clk, r2592_out, r2593_out);
	reg32 r2594 (rst, clk, r2593_out, r2594_out);
	reg32 r2595 (rst, clk, r2594_out, r2595_out);
	reg32 r2596 (rst, clk, r2595_out, r2596_out);
	reg32 r2597 (rst, clk, r2596_out, r2597_out);
	reg32 r2598 (rst, clk, r2597_out, r2598_out);
	reg32 r2599 (rst, clk, r2598_out, r2599_out);
	reg32 r2600 (rst, clk, r2599_out, r2600_out);
	reg32 r2601 (rst, clk, r2600_out, r2601_out);
	reg32 r2602 (rst, clk, r2601_out, r2602_out);
	reg32 r2603 (rst, clk, r2602_out, r2603_out);
	reg32 r2604 (rst, clk, r2603_out, r2604_out);
	reg32 r2605 (rst, clk, r2604_out, r2605_out);
	reg32 r2606 (rst, clk, r2605_out, r2606_out);
	reg32 r2607 (rst, clk, r2606_out, r2607_out);
	reg32 r2608 (rst, clk, r2607_out, r2608_out);
	reg32 r2609 (rst, clk, r2608_out, r2609_out);
	reg32 r2610 (rst, clk, r2609_out, r2610_out);
	reg32 r2611 (rst, clk, r2610_out, r2611_out);
	reg32 r2612 (rst, clk, r2611_out, r2612_out);
	reg32 r2613 (rst, clk, r2612_out, r2613_out);
	reg32 r2614 (rst, clk, r2613_out, r2614_out);
	reg32 r2615 (rst, clk, r2614_out, r2615_out);
	reg32 r2616 (rst, clk, r2615_out, r2616_out);
	reg32 r2617 (rst, clk, r2616_out, r2617_out);
	reg32 r2618 (rst, clk, r2617_out, r2618_out);
	reg32 r2619 (rst, clk, r2618_out, r2619_out);
	reg32 r2620 (rst, clk, r2619_out, r2620_out);
	reg32 r2621 (rst, clk, r2620_out, r2621_out);
	reg32 r2622 (rst, clk, r2621_out, r2622_out);
	reg32 r2623 (rst, clk, r2622_out, r2623_out);
	reg32 r2624 (rst, clk, r2623_out, r2624_out);
	reg32 r2625 (rst, clk, r2624_out, r2625_out);
	reg32 r2626 (rst, clk, r2625_out, r2626_out);
	reg32 r2627 (rst, clk, r2626_out, r2627_out);
	reg32 r2628 (rst, clk, r2627_out, r2628_out);
	reg32 r2629 (rst, clk, r2628_out, r2629_out);
	reg32 r2630 (rst, clk, r2629_out, r2630_out);
	reg32 r2631 (rst, clk, r2630_out, r2631_out);
	reg32 r2632 (rst, clk, r2631_out, r2632_out);
	reg32 r2633 (rst, clk, r2632_out, r2633_out);
	reg32 r2634 (rst, clk, r2633_out, r2634_out);
	reg32 r2635 (rst, clk, r2634_out, r2635_out);
	reg32 r2636 (rst, clk, r2635_out, r2636_out);
	reg32 r2637 (rst, clk, r2636_out, r2637_out);
	reg32 r2638 (rst, clk, r2637_out, r2638_out);
	reg32 r2639 (rst, clk, r2638_out, r2639_out);
	reg32 r2640 (rst, clk, r2639_out, r2640_out);
	reg32 r2641 (rst, clk, r2640_out, r2641_out);
	reg32 r2642 (rst, clk, r2641_out, r2642_out);
	reg32 r2643 (rst, clk, r2642_out, r2643_out);
	reg32 r2644 (rst, clk, r2643_out, r2644_out);
	reg32 r2645 (rst, clk, r2644_out, r2645_out);
	reg32 r2646 (rst, clk, r2645_out, r2646_out);
	reg32 r2647 (rst, clk, r2646_out, r2647_out);
	reg32 r2648 (rst, clk, r2647_out, r2648_out);
	reg32 r2649 (rst, clk, r2648_out, r2649_out);
	reg32 r2650 (rst, clk, r2649_out, r2650_out);
	reg32 r2651 (rst, clk, r2650_out, r2651_out);
	reg32 r2652 (rst, clk, r2651_out, r2652_out);
	reg32 r2653 (rst, clk, r2652_out, r2653_out);
	reg32 r2654 (rst, clk, r2653_out, r2654_out);
	reg32 r2655 (rst, clk, r2654_out, r2655_out);
	reg32 r2656 (rst, clk, r2655_out, r2656_out);
	reg32 r2657 (rst, clk, r2656_out, r2657_out);
	reg32 r2658 (rst, clk, r2657_out, r2658_out);
	reg32 r2659 (rst, clk, r2658_out, r2659_out);
	reg32 r2660 (rst, clk, r2659_out, r2660_out);
	reg32 r2661 (rst, clk, r2660_out, r2661_out);
	reg32 r2662 (rst, clk, r2661_out, r2662_out);
	reg32 r2663 (rst, clk, r2662_out, r2663_out);
	reg32 r2664 (rst, clk, r2663_out, r2664_out);
	reg32 r2665 (rst, clk, r2664_out, r2665_out);
	reg32 r2666 (rst, clk, r2665_out, r2666_out);
	reg32 r2667 (rst, clk, r2666_out, r2667_out);
	reg32 r2668 (rst, clk, r2667_out, r2668_out);
	reg32 r2669 (rst, clk, r2668_out, r2669_out);
	reg32 r2670 (rst, clk, r2669_out, r2670_out);
	reg32 r2671 (rst, clk, r2670_out, r2671_out);
	reg32 r2672 (rst, clk, r2671_out, r2672_out);
	reg32 r2673 (rst, clk, r2672_out, r2673_out);
	reg32 r2674 (rst, clk, r2673_out, r2674_out);
	reg32 r2675 (rst, clk, r2674_out, r2675_out);
	reg32 r2676 (rst, clk, r2675_out, r2676_out);
	reg32 r2677 (rst, clk, r2676_out, r2677_out);
	reg32 r2678 (rst, clk, r2677_out, r2678_out);
	reg32 r2679 (rst, clk, r2678_out, r2679_out);
	reg32 r2680 (rst, clk, r2679_out, r2680_out);
	reg32 r2681 (rst, clk, r2680_out, r2681_out);
	reg32 r2682 (rst, clk, r2681_out, r2682_out);
	reg32 r2683 (rst, clk, r2682_out, r2683_out);
	reg32 r2684 (rst, clk, r2683_out, r2684_out);
	reg32 r2685 (rst, clk, r2684_out, r2685_out);
	reg32 r2686 (rst, clk, r2685_out, r2686_out);
	reg32 r2687 (rst, clk, r2686_out, r2687_out);
	reg32 r2688 (rst, clk, r2687_out, r2688_out);
	reg32 r2689 (rst, clk, r2688_out, r2689_out);
	reg32 r2690 (rst, clk, r2689_out, r2690_out);
	reg32 r2691 (rst, clk, r2690_out, r2691_out);
	reg32 r2692 (rst, clk, r2691_out, r2692_out);
	reg32 r2693 (rst, clk, r2692_out, r2693_out);
	reg32 r2694 (rst, clk, r2693_out, r2694_out);
	reg32 r2695 (rst, clk, r2694_out, r2695_out);
	reg32 r2696 (rst, clk, r2695_out, r2696_out);
	reg32 r2697 (rst, clk, r2696_out, r2697_out);
	reg32 r2698 (rst, clk, r2697_out, r2698_out);
	reg32 r2699 (rst, clk, r2698_out, r2699_out);
	reg32 r2700 (rst, clk, r2699_out, r2700_out);
	reg32 r2701 (rst, clk, r2700_out, r2701_out);
	reg32 r2702 (rst, clk, r2701_out, r2702_out);
	reg32 r2703 (rst, clk, r2702_out, r2703_out);
	reg32 r2704 (rst, clk, r2703_out, r2704_out);
	reg32 r2705 (rst, clk, r2704_out, r2705_out);
	reg32 r2706 (rst, clk, r2705_out, r2706_out);
	reg32 r2707 (rst, clk, r2706_out, r2707_out);
	reg32 r2708 (rst, clk, r2707_out, r2708_out);
	reg32 r2709 (rst, clk, r2708_out, r2709_out);
	reg32 r2710 (rst, clk, r2709_out, r2710_out);
	reg32 r2711 (rst, clk, r2710_out, r2711_out);
	reg32 r2712 (rst, clk, r2711_out, r2712_out);
	reg32 r2713 (rst, clk, r2712_out, r2713_out);
	reg32 r2714 (rst, clk, r2713_out, r2714_out);
	reg32 r2715 (rst, clk, r2714_out, r2715_out);
	reg32 r2716 (rst, clk, r2715_out, r2716_out);
	reg32 r2717 (rst, clk, r2716_out, r2717_out);
	reg32 r2718 (rst, clk, r2717_out, r2718_out);
	reg32 r2719 (rst, clk, r2718_out, r2719_out);
	reg32 r2720 (rst, clk, r2719_out, r2720_out);
	reg32 r2721 (rst, clk, r2720_out, r2721_out);
	reg32 r2722 (rst, clk, r2721_out, r2722_out);
	reg32 r2723 (rst, clk, r2722_out, r2723_out);
	reg32 r2724 (rst, clk, r2723_out, r2724_out);
	reg32 r2725 (rst, clk, r2724_out, r2725_out);
	reg32 r2726 (rst, clk, r2725_out, r2726_out);
	reg32 r2727 (rst, clk, r2726_out, r2727_out);
	reg32 r2728 (rst, clk, r2727_out, r2728_out);
	reg32 r2729 (rst, clk, r2728_out, r2729_out);
	reg32 r2730 (rst, clk, r2729_out, r2730_out);
	reg32 r2731 (rst, clk, r2730_out, r2731_out);
	reg32 r2732 (rst, clk, r2731_out, r2732_out);
	reg32 r2733 (rst, clk, r2732_out, r2733_out);
	reg32 r2734 (rst, clk, r2733_out, r2734_out);
	reg32 r2735 (rst, clk, r2734_out, r2735_out);
	reg32 r2736 (rst, clk, r2735_out, r2736_out);
	reg32 r2737 (rst, clk, r2736_out, r2737_out);
	reg32 r2738 (rst, clk, r2737_out, r2738_out);
	reg32 r2739 (rst, clk, r2738_out, r2739_out);
	reg32 r2740 (rst, clk, r2739_out, r2740_out);
	reg32 r2741 (rst, clk, r2740_out, r2741_out);
	reg32 r2742 (rst, clk, r2741_out, r2742_out);
	reg32 r2743 (rst, clk, r2742_out, r2743_out);
	reg32 r2744 (rst, clk, r2743_out, r2744_out);
	reg32 r2745 (rst, clk, r2744_out, r2745_out);
	reg32 r2746 (rst, clk, r2745_out, r2746_out);
	reg32 r2747 (rst, clk, r2746_out, r2747_out);
	reg32 r2748 (rst, clk, r2747_out, r2748_out);
	reg32 r2749 (rst, clk, r2748_out, r2749_out);
	reg32 r2750 (rst, clk, r2749_out, r2750_out);
	reg32 r2751 (rst, clk, r2750_out, r2751_out);
	reg32 r2752 (rst, clk, r2751_out, r2752_out);
	reg32 r2753 (rst, clk, r2752_out, r2753_out);
	reg32 r2754 (rst, clk, r2753_out, r2754_out);
	reg32 r2755 (rst, clk, r2754_out, r2755_out);
	reg32 r2756 (rst, clk, r2755_out, r2756_out);
	reg32 r2757 (rst, clk, r2756_out, r2757_out);
	reg32 r2758 (rst, clk, r2757_out, r2758_out);
	reg32 r2759 (rst, clk, r2758_out, r2759_out);
	reg32 r2760 (rst, clk, r2759_out, r2760_out);
	reg32 r2761 (rst, clk, r2760_out, r2761_out);
	reg32 r2762 (rst, clk, r2761_out, r2762_out);
	reg32 r2763 (rst, clk, r2762_out, r2763_out);
	reg32 r2764 (rst, clk, r2763_out, r2764_out);
	reg32 r2765 (rst, clk, r2764_out, r2765_out);
	reg32 r2766 (rst, clk, r2765_out, r2766_out);
	reg32 r2767 (rst, clk, r2766_out, r2767_out);
	reg32 r2768 (rst, clk, r2767_out, r2768_out);
	reg32 r2769 (rst, clk, r2768_out, r2769_out);
	reg32 r2770 (rst, clk, r2769_out, r2770_out);
	reg32 r2771 (rst, clk, r2770_out, r2771_out);
	reg32 r2772 (rst, clk, r2771_out, r2772_out);
	reg32 r2773 (rst, clk, r2772_out, r2773_out);
	reg32 r2774 (rst, clk, r2773_out, r2774_out);
	reg32 r2775 (rst, clk, r2774_out, r2775_out);
	reg32 r2776 (rst, clk, r2775_out, r2776_out);
	reg32 r2777 (rst, clk, r2776_out, r2777_out);
	reg32 r2778 (rst, clk, r2777_out, r2778_out);
	reg32 r2779 (rst, clk, r2778_out, r2779_out);
	reg32 r2780 (rst, clk, r2779_out, r2780_out);
	reg32 r2781 (rst, clk, r2780_out, r2781_out);
	reg32 r2782 (rst, clk, r2781_out, r2782_out);
	reg32 r2783 (rst, clk, r2782_out, r2783_out);
	reg32 r2784 (rst, clk, r2783_out, r2784_out);
	reg32 r2785 (rst, clk, r2784_out, r2785_out);
	reg32 r2786 (rst, clk, r2785_out, r2786_out);
	reg32 r2787 (rst, clk, r2786_out, r2787_out);
	reg32 r2788 (rst, clk, r2787_out, r2788_out);
	reg32 r2789 (rst, clk, r2788_out, r2789_out);
	reg32 r2790 (rst, clk, r2789_out, r2790_out);
	reg32 r2791 (rst, clk, r2790_out, r2791_out);
	reg32 r2792 (rst, clk, r2791_out, r2792_out);
	reg32 r2793 (rst, clk, r2792_out, r2793_out);
	reg32 r2794 (rst, clk, r2793_out, r2794_out);
	reg32 r2795 (rst, clk, r2794_out, r2795_out);
	reg32 r2796 (rst, clk, r2795_out, r2796_out);
	reg32 r2797 (rst, clk, r2796_out, r2797_out);
	reg32 r2798 (rst, clk, r2797_out, r2798_out);
	reg32 r2799 (rst, clk, r2798_out, r2799_out);
	reg32 r2800 (rst, clk, r2799_out, r2800_out);
	reg32 r2801 (rst, clk, r2800_out, r2801_out);
	reg32 r2802 (rst, clk, r2801_out, r2802_out);
	reg32 r2803 (rst, clk, r2802_out, r2803_out);
	reg32 r2804 (rst, clk, r2803_out, r2804_out);
	reg32 r2805 (rst, clk, r2804_out, r2805_out);
	reg32 r2806 (rst, clk, r2805_out, r2806_out);
	reg32 r2807 (rst, clk, r2806_out, r2807_out);
	reg32 r2808 (rst, clk, r2807_out, r2808_out);
	reg32 r2809 (rst, clk, r2808_out, r2809_out);
	reg32 r2810 (rst, clk, r2809_out, r2810_out);
	reg32 r2811 (rst, clk, r2810_out, r2811_out);
	reg32 r2812 (rst, clk, r2811_out, r2812_out);
	reg32 r2813 (rst, clk, r2812_out, r2813_out);
	reg32 r2814 (rst, clk, r2813_out, r2814_out);
	reg32 r2815 (rst, clk, r2814_out, r2815_out);
	reg32 r2816 (rst, clk, r2815_out, r2816_out);
	reg32 r2817 (rst, clk, r2816_out, r2817_out);
	reg32 r2818 (rst, clk, r2817_out, r2818_out);
	reg32 r2819 (rst, clk, r2818_out, r2819_out);
	reg32 r2820 (rst, clk, r2819_out, r2820_out);
	reg32 r2821 (rst, clk, r2820_out, r2821_out);
	reg32 r2822 (rst, clk, r2821_out, r2822_out);
	reg32 r2823 (rst, clk, r2822_out, r2823_out);
	reg32 r2824 (rst, clk, r2823_out, r2824_out);
	reg32 r2825 (rst, clk, r2824_out, r2825_out);
	reg32 r2826 (rst, clk, r2825_out, r2826_out);
	reg32 r2827 (rst, clk, r2826_out, r2827_out);
	reg32 r2828 (rst, clk, r2827_out, r2828_out);
	reg32 r2829 (rst, clk, r2828_out, r2829_out);
	reg32 r2830 (rst, clk, r2829_out, r2830_out);
	reg32 r2831 (rst, clk, r2830_out, r2831_out);
	reg32 r2832 (rst, clk, r2831_out, r2832_out);
	reg32 r2833 (rst, clk, r2832_out, r2833_out);
	reg32 r2834 (rst, clk, r2833_out, r2834_out);
	reg32 r2835 (rst, clk, r2834_out, r2835_out);
	reg32 r2836 (rst, clk, r2835_out, r2836_out);
	reg32 r2837 (rst, clk, r2836_out, r2837_out);
	reg32 r2838 (rst, clk, r2837_out, r2838_out);
	reg32 r2839 (rst, clk, r2838_out, r2839_out);
	reg32 r2840 (rst, clk, r2839_out, r2840_out);
	reg32 r2841 (rst, clk, r2840_out, r2841_out);
	reg32 r2842 (rst, clk, r2841_out, r2842_out);
	reg32 r2843 (rst, clk, r2842_out, r2843_out);
	reg32 r2844 (rst, clk, r2843_out, r2844_out);
	reg32 r2845 (rst, clk, r2844_out, r2845_out);
	reg32 r2846 (rst, clk, r2845_out, r2846_out);
	reg32 r2847 (rst, clk, r2846_out, r2847_out);
	reg32 r2848 (rst, clk, r2847_out, r2848_out);
	reg32 r2849 (rst, clk, r2848_out, r2849_out);
	reg32 r2850 (rst, clk, r2849_out, r2850_out);
	reg32 r2851 (rst, clk, r2850_out, r2851_out);
	reg32 r2852 (rst, clk, r2851_out, r2852_out);
	reg32 r2853 (rst, clk, r2852_out, r2853_out);
	reg32 r2854 (rst, clk, r2853_out, r2854_out);
	reg32 r2855 (rst, clk, r2854_out, r2855_out);
	reg32 r2856 (rst, clk, r2855_out, r2856_out);
	reg32 r2857 (rst, clk, r2856_out, r2857_out);
	reg32 r2858 (rst, clk, r2857_out, r2858_out);
	reg32 r2859 (rst, clk, r2858_out, r2859_out);
	reg32 r2860 (rst, clk, r2859_out, r2860_out);
	reg32 r2861 (rst, clk, r2860_out, r2861_out);
	reg32 r2862 (rst, clk, r2861_out, r2862_out);
	reg32 r2863 (rst, clk, r2862_out, r2863_out);
	reg32 r2864 (rst, clk, r2863_out, r2864_out);
	reg32 r2865 (rst, clk, r2864_out, r2865_out);
	reg32 r2866 (rst, clk, r2865_out, r2866_out);
	reg32 r2867 (rst, clk, r2866_out, r2867_out);
	reg32 r2868 (rst, clk, r2867_out, r2868_out);
	reg32 r2869 (rst, clk, r2868_out, r2869_out);
	reg32 r2870 (rst, clk, r2869_out, r2870_out);
	reg32 r2871 (rst, clk, r2870_out, r2871_out);
	reg32 r2872 (rst, clk, r2871_out, r2872_out);
	reg32 r2873 (rst, clk, r2872_out, r2873_out);
	reg32 r2874 (rst, clk, r2873_out, r2874_out);
	reg32 r2875 (rst, clk, r2874_out, r2875_out);
	reg32 r2876 (rst, clk, r2875_out, r2876_out);
	reg32 r2877 (rst, clk, r2876_out, r2877_out);
	reg32 r2878 (rst, clk, r2877_out, r2878_out);
	reg32 r2879 (rst, clk, r2878_out, r2879_out);
	reg32 r2880 (rst, clk, r2879_out, r2880_out);
	reg32 r2881 (rst, clk, r2880_out, r2881_out);
	reg32 r2882 (rst, clk, r2881_out, r2882_out);
	reg32 r2883 (rst, clk, r2882_out, r2883_out);
	reg32 r2884 (rst, clk, r2883_out, r2884_out);
	reg32 r2885 (rst, clk, r2884_out, r2885_out);
	reg32 r2886 (rst, clk, r2885_out, r2886_out);
	reg32 r2887 (rst, clk, r2886_out, r2887_out);
	reg32 r2888 (rst, clk, r2887_out, r2888_out);
	reg32 r2889 (rst, clk, r2888_out, r2889_out);
	reg32 r2890 (rst, clk, r2889_out, r2890_out);
	reg32 r2891 (rst, clk, r2890_out, r2891_out);
	reg32 r2892 (rst, clk, r2891_out, r2892_out);
	reg32 r2893 (rst, clk, r2892_out, r2893_out);
	reg32 r2894 (rst, clk, r2893_out, r2894_out);
	reg32 r2895 (rst, clk, r2894_out, r2895_out);
	reg32 r2896 (rst, clk, r2895_out, r2896_out);
	reg32 r2897 (rst, clk, r2896_out, r2897_out);
	reg32 r2898 (rst, clk, r2897_out, r2898_out);
	reg32 r2899 (rst, clk, r2898_out, r2899_out);
	reg32 r2900 (rst, clk, r2899_out, r2900_out);
	reg32 r2901 (rst, clk, r2900_out, r2901_out);
	reg32 r2902 (rst, clk, r2901_out, r2902_out);
	reg32 r2903 (rst, clk, r2902_out, r2903_out);
	reg32 r2904 (rst, clk, r2903_out, r2904_out);
	reg32 r2905 (rst, clk, r2904_out, r2905_out);
	reg32 r2906 (rst, clk, r2905_out, r2906_out);
	reg32 r2907 (rst, clk, r2906_out, r2907_out);
	reg32 r2908 (rst, clk, r2907_out, r2908_out);
	reg32 r2909 (rst, clk, r2908_out, r2909_out);
	reg32 r2910 (rst, clk, r2909_out, r2910_out);
	reg32 r2911 (rst, clk, r2910_out, r2911_out);
	reg32 r2912 (rst, clk, r2911_out, r2912_out);
	reg32 r2913 (rst, clk, r2912_out, r2913_out);
	reg32 r2914 (rst, clk, r2913_out, r2914_out);
	reg32 r2915 (rst, clk, r2914_out, r2915_out);
	reg32 r2916 (rst, clk, r2915_out, r2916_out);
	reg32 r2917 (rst, clk, r2916_out, r2917_out);
	reg32 r2918 (rst, clk, r2917_out, r2918_out);
	reg32 r2919 (rst, clk, r2918_out, r2919_out);
	reg32 r2920 (rst, clk, r2919_out, r2920_out);
	reg32 r2921 (rst, clk, r2920_out, r2921_out);
	reg32 r2922 (rst, clk, r2921_out, r2922_out);
	reg32 r2923 (rst, clk, r2922_out, r2923_out);
	reg32 r2924 (rst, clk, r2923_out, r2924_out);
	reg32 r2925 (rst, clk, r2924_out, r2925_out);
	reg32 r2926 (rst, clk, r2925_out, r2926_out);
	reg32 r2927 (rst, clk, r2926_out, r2927_out);
	reg32 r2928 (rst, clk, r2927_out, r2928_out);
	reg32 r2929 (rst, clk, r2928_out, r2929_out);
	reg32 r2930 (rst, clk, r2929_out, r2930_out);
	reg32 r2931 (rst, clk, r2930_out, r2931_out);
	reg32 r2932 (rst, clk, r2931_out, r2932_out);
	reg32 r2933 (rst, clk, r2932_out, r2933_out);
	reg32 r2934 (rst, clk, r2933_out, r2934_out);
	reg32 r2935 (rst, clk, r2934_out, r2935_out);
	reg32 r2936 (rst, clk, r2935_out, r2936_out);
	reg32 r2937 (rst, clk, r2936_out, r2937_out);
	reg32 r2938 (rst, clk, r2937_out, r2938_out);
	reg32 r2939 (rst, clk, r2938_out, r2939_out);
	reg32 r2940 (rst, clk, r2939_out, r2940_out);
	reg32 r2941 (rst, clk, r2940_out, r2941_out);
	reg32 r2942 (rst, clk, r2941_out, r2942_out);
	reg32 r2943 (rst, clk, r2942_out, r2943_out);
	reg32 r2944 (rst, clk, r2943_out, r2944_out);
	reg32 r2945 (rst, clk, r2944_out, r2945_out);
	reg32 r2946 (rst, clk, r2945_out, r2946_out);
	reg32 r2947 (rst, clk, r2946_out, r2947_out);
	reg32 r2948 (rst, clk, r2947_out, r2948_out);
	reg32 r2949 (rst, clk, r2948_out, r2949_out);
	reg32 r2950 (rst, clk, r2949_out, r2950_out);
	reg32 r2951 (rst, clk, r2950_out, r2951_out);
	reg32 r2952 (rst, clk, r2951_out, r2952_out);
	reg32 r2953 (rst, clk, r2952_out, r2953_out);
	reg32 r2954 (rst, clk, r2953_out, r2954_out);
	reg32 r2955 (rst, clk, r2954_out, r2955_out);
	reg32 r2956 (rst, clk, r2955_out, r2956_out);
	reg32 r2957 (rst, clk, r2956_out, r2957_out);
	reg32 r2958 (rst, clk, r2957_out, r2958_out);
	reg32 r2959 (rst, clk, r2958_out, r2959_out);
	reg32 r2960 (rst, clk, r2959_out, r2960_out);
	reg32 r2961 (rst, clk, r2960_out, r2961_out);
	reg32 r2962 (rst, clk, r2961_out, r2962_out);
	reg32 r2963 (rst, clk, r2962_out, r2963_out);
	reg32 r2964 (rst, clk, r2963_out, r2964_out);
	reg32 r2965 (rst, clk, r2964_out, r2965_out);
	reg32 r2966 (rst, clk, r2965_out, r2966_out);
	reg32 r2967 (rst, clk, r2966_out, r2967_out);
	reg32 r2968 (rst, clk, r2967_out, r2968_out);
	reg32 r2969 (rst, clk, r2968_out, r2969_out);
	reg32 r2970 (rst, clk, r2969_out, r2970_out);
	reg32 r2971 (rst, clk, r2970_out, r2971_out);
	reg32 r2972 (rst, clk, r2971_out, r2972_out);
	reg32 r2973 (rst, clk, r2972_out, r2973_out);
	reg32 r2974 (rst, clk, r2973_out, r2974_out);
	reg32 r2975 (rst, clk, r2974_out, r2975_out);
	reg32 r2976 (rst, clk, r2975_out, r2976_out);
	reg32 r2977 (rst, clk, r2976_out, r2977_out);
	reg32 r2978 (rst, clk, r2977_out, r2978_out);
	reg32 r2979 (rst, clk, r2978_out, r2979_out);
	reg32 r2980 (rst, clk, r2979_out, r2980_out);
	reg32 r2981 (rst, clk, r2980_out, r2981_out);
	reg32 r2982 (rst, clk, r2981_out, r2982_out);
	reg32 r2983 (rst, clk, r2982_out, r2983_out);
	reg32 r2984 (rst, clk, r2983_out, r2984_out);
	reg32 r2985 (rst, clk, r2984_out, r2985_out);
	reg32 r2986 (rst, clk, r2985_out, r2986_out);
	reg32 r2987 (rst, clk, r2986_out, r2987_out);
	reg32 r2988 (rst, clk, r2987_out, r2988_out);
	reg32 r2989 (rst, clk, r2988_out, r2989_out);
	reg32 r2990 (rst, clk, r2989_out, r2990_out);
	reg32 r2991 (rst, clk, r2990_out, r2991_out);
	reg32 r2992 (rst, clk, r2991_out, r2992_out);
	reg32 r2993 (rst, clk, r2992_out, r2993_out);
	reg32 r2994 (rst, clk, r2993_out, r2994_out);
	reg32 r2995 (rst, clk, r2994_out, r2995_out);
	reg32 r2996 (rst, clk, r2995_out, r2996_out);
	reg32 r2997 (rst, clk, r2996_out, r2997_out);
	reg32 r2998 (rst, clk, r2997_out, r2998_out);
	reg32 r2999 (rst, clk, r2998_out, r2999_out);

	assign out = r2999_out;
endmodule
