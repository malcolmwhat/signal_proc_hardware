module reg100 ( in, clk, rst, out );
	input[31:0] in;
	input clk;
	input rst;
	output[31:0] out;

	wire [31:0] r0_out;
	wire [31:0] r1_out;
	wire [31:0] r2_out;
	wire [31:0] r3_out;
	wire [31:0] r4_out;
	wire [31:0] r5_out;
	wire [31:0] r6_out;
	wire [31:0] r7_out;
	wire [31:0] r8_out;
	wire [31:0] r9_out;
	wire [31:0] r10_out;
	wire [31:0] r11_out;
	wire [31:0] r12_out;
	wire [31:0] r13_out;
	wire [31:0] r14_out;
	wire [31:0] r15_out;
	wire [31:0] r16_out;
	wire [31:0] r17_out;
	wire [31:0] r18_out;
	wire [31:0] r19_out;
	wire [31:0] r20_out;
	wire [31:0] r21_out;
	wire [31:0] r22_out;
	wire [31:0] r23_out;
	wire [31:0] r24_out;
	wire [31:0] r25_out;
	wire [31:0] r26_out;
	wire [31:0] r27_out;
	wire [31:0] r28_out;
	wire [31:0] r29_out;
	wire [31:0] r30_out;
	wire [31:0] r31_out;
	wire [31:0] r32_out;
	wire [31:0] r33_out;
	wire [31:0] r34_out;
	wire [31:0] r35_out;
	wire [31:0] r36_out;
	wire [31:0] r37_out;
	wire [31:0] r38_out;
	wire [31:0] r39_out;
	wire [31:0] r40_out;
	wire [31:0] r41_out;
	wire [31:0] r42_out;
	wire [31:0] r43_out;
	wire [31:0] r44_out;
	wire [31:0] r45_out;
	wire [31:0] r46_out;
	wire [31:0] r47_out;
	wire [31:0] r48_out;
	wire [31:0] r49_out;
	wire [31:0] r50_out;
	wire [31:0] r51_out;
	wire [31:0] r52_out;
	wire [31:0] r53_out;
	wire [31:0] r54_out;
	wire [31:0] r55_out;
	wire [31:0] r56_out;
	wire [31:0] r57_out;
	wire [31:0] r58_out;
	wire [31:0] r59_out;
	wire [31:0] r60_out;
	wire [31:0] r61_out;
	wire [31:0] r62_out;
	wire [31:0] r63_out;
	wire [31:0] r64_out;
	wire [31:0] r65_out;
	wire [31:0] r66_out;
	wire [31:0] r67_out;
	wire [31:0] r68_out;
	wire [31:0] r69_out;
	wire [31:0] r70_out;
	wire [31:0] r71_out;
	wire [31:0] r72_out;
	wire [31:0] r73_out;
	wire [31:0] r74_out;
	wire [31:0] r75_out;
	wire [31:0] r76_out;
	wire [31:0] r77_out;
	wire [31:0] r78_out;
	wire [31:0] r79_out;
	wire [31:0] r80_out;
	wire [31:0] r81_out;
	wire [31:0] r82_out;
	wire [31:0] r83_out;
	wire [31:0] r84_out;
	wire [31:0] r85_out;
	wire [31:0] r86_out;
	wire [31:0] r87_out;
	wire [31:0] r88_out;
	wire [31:0] r89_out;
	wire [31:0] r90_out;
	wire [31:0] r91_out;
	wire [31:0] r92_out;
	wire [31:0] r93_out;
	wire [31:0] r94_out;
	wire [31:0] r95_out;
	wire [31:0] r96_out;
	wire [31:0] r97_out;
	wire [31:0] r98_out;
	wire [31:0] r99_out;

	reg32 r0 (rst, clk, in, r0_out);
	reg32 r1 (rst, clk, r0_out, r1_out);
	reg32 r2 (rst, clk, r1_out, r2_out);
	reg32 r3 (rst, clk, r2_out, r3_out);
	reg32 r4 (rst, clk, r3_out, r4_out);
	reg32 r5 (rst, clk, r4_out, r5_out);
	reg32 r6 (rst, clk, r5_out, r6_out);
	reg32 r7 (rst, clk, r6_out, r7_out);
	reg32 r8 (rst, clk, r7_out, r8_out);
	reg32 r9 (rst, clk, r8_out, r9_out);
	reg32 r10 (rst, clk, r9_out, r10_out);
	reg32 r11 (rst, clk, r10_out, r11_out);
	reg32 r12 (rst, clk, r11_out, r12_out);
	reg32 r13 (rst, clk, r12_out, r13_out);
	reg32 r14 (rst, clk, r13_out, r14_out);
	reg32 r15 (rst, clk, r14_out, r15_out);
	reg32 r16 (rst, clk, r15_out, r16_out);
	reg32 r17 (rst, clk, r16_out, r17_out);
	reg32 r18 (rst, clk, r17_out, r18_out);
	reg32 r19 (rst, clk, r18_out, r19_out);
	reg32 r20 (rst, clk, r19_out, r20_out);
	reg32 r21 (rst, clk, r20_out, r21_out);
	reg32 r22 (rst, clk, r21_out, r22_out);
	reg32 r23 (rst, clk, r22_out, r23_out);
	reg32 r24 (rst, clk, r23_out, r24_out);
	reg32 r25 (rst, clk, r24_out, r25_out);
	reg32 r26 (rst, clk, r25_out, r26_out);
	reg32 r27 (rst, clk, r26_out, r27_out);
	reg32 r28 (rst, clk, r27_out, r28_out);
	reg32 r29 (rst, clk, r28_out, r29_out);
	reg32 r30 (rst, clk, r29_out, r30_out);
	reg32 r31 (rst, clk, r30_out, r31_out);
	reg32 r32 (rst, clk, r31_out, r32_out);
	reg32 r33 (rst, clk, r32_out, r33_out);
	reg32 r34 (rst, clk, r33_out, r34_out);
	reg32 r35 (rst, clk, r34_out, r35_out);
	reg32 r36 (rst, clk, r35_out, r36_out);
	reg32 r37 (rst, clk, r36_out, r37_out);
	reg32 r38 (rst, clk, r37_out, r38_out);
	reg32 r39 (rst, clk, r38_out, r39_out);
	reg32 r40 (rst, clk, r39_out, r40_out);
	reg32 r41 (rst, clk, r40_out, r41_out);
	reg32 r42 (rst, clk, r41_out, r42_out);
	reg32 r43 (rst, clk, r42_out, r43_out);
	reg32 r44 (rst, clk, r43_out, r44_out);
	reg32 r45 (rst, clk, r44_out, r45_out);
	reg32 r46 (rst, clk, r45_out, r46_out);
	reg32 r47 (rst, clk, r46_out, r47_out);
	reg32 r48 (rst, clk, r47_out, r48_out);
	reg32 r49 (rst, clk, r48_out, r49_out);
	reg32 r50 (rst, clk, r49_out, r50_out);
	reg32 r51 (rst, clk, r50_out, r51_out);
	reg32 r52 (rst, clk, r51_out, r52_out);
	reg32 r53 (rst, clk, r52_out, r53_out);
	reg32 r54 (rst, clk, r53_out, r54_out);
	reg32 r55 (rst, clk, r54_out, r55_out);
	reg32 r56 (rst, clk, r55_out, r56_out);
	reg32 r57 (rst, clk, r56_out, r57_out);
	reg32 r58 (rst, clk, r57_out, r58_out);
	reg32 r59 (rst, clk, r58_out, r59_out);
	reg32 r60 (rst, clk, r59_out, r60_out);
	reg32 r61 (rst, clk, r60_out, r61_out);
	reg32 r62 (rst, clk, r61_out, r62_out);
	reg32 r63 (rst, clk, r62_out, r63_out);
	reg32 r64 (rst, clk, r63_out, r64_out);
	reg32 r65 (rst, clk, r64_out, r65_out);
	reg32 r66 (rst, clk, r65_out, r66_out);
	reg32 r67 (rst, clk, r66_out, r67_out);
	reg32 r68 (rst, clk, r67_out, r68_out);
	reg32 r69 (rst, clk, r68_out, r69_out);
	reg32 r70 (rst, clk, r69_out, r70_out);
	reg32 r71 (rst, clk, r70_out, r71_out);
	reg32 r72 (rst, clk, r71_out, r72_out);
	reg32 r73 (rst, clk, r72_out, r73_out);
	reg32 r74 (rst, clk, r73_out, r74_out);
	reg32 r75 (rst, clk, r74_out, r75_out);
	reg32 r76 (rst, clk, r75_out, r76_out);
	reg32 r77 (rst, clk, r76_out, r77_out);
	reg32 r78 (rst, clk, r77_out, r78_out);
	reg32 r79 (rst, clk, r78_out, r79_out);
	reg32 r80 (rst, clk, r79_out, r80_out);
	reg32 r81 (rst, clk, r80_out, r81_out);
	reg32 r82 (rst, clk, r81_out, r82_out);
	reg32 r83 (rst, clk, r82_out, r83_out);
	reg32 r84 (rst, clk, r83_out, r84_out);
	reg32 r85 (rst, clk, r84_out, r85_out);
	reg32 r86 (rst, clk, r85_out, r86_out);
	reg32 r87 (rst, clk, r86_out, r87_out);
	reg32 r88 (rst, clk, r87_out, r88_out);
	reg32 r89 (rst, clk, r88_out, r89_out);
	reg32 r90 (rst, clk, r89_out, r90_out);
	reg32 r91 (rst, clk, r90_out, r91_out);
	reg32 r92 (rst, clk, r91_out, r92_out);
	reg32 r93 (rst, clk, r92_out, r93_out);
	reg32 r94 (rst, clk, r93_out, r94_out);
	reg32 r95 (rst, clk, r94_out, r95_out);
	reg32 r96 (rst, clk, r95_out, r96_out);
	reg32 r97 (rst, clk, r96_out, r97_out);
	reg32 r98 (rst, clk, r97_out, r98_out);
	reg32 r99 (rst, clk, r98_out, r99_out);

	assign out = r99_out;
endmodule
